
module alu ( a, b, op, result, zero );
  input [31:0] a;
  input [31:0] b;
  input [3:0] op;
  output [31:0] result;
  output zero;
  wire   n7897, sel, n509, n3158, net211934, net211935, net211939, net211942,
         net211946, net211949, net211950, net211993, net211994, net212005,
         net212007, net212008, net212010, net212023, net212061, net212092,
         net212093, net212094, net212102, net212114, net212116, net212121,
         net212125, net212126, net212128, net212129, net212134, net212137,
         net212138, net212140, net212141, net212143, net212145, net212146,
         net212283, net212284, net212377, net212381, net212383, net212391,
         net212392, net212393, net212394, net212411, net212412, net212420,
         net212433, net212437, net212438, net212442, net212443, net212447,
         net212448, net212451, net212468, net212470, net212483, net212485,
         net212493, net212495, net212634, net212635, net212636, net212645,
         net212646, net212649, net212651, net212652, net212653, net212655,
         net212656, net212660, net212672, net212673, net212674, net212677,
         net212679, net212681, net212685, net212686, net212688, net212689,
         net212690, net212691, net212693, net212694, net212696, net212697,
         net212698, net212700, net212703, net212704, net212705, net212735,
         net212738, net212739, net212740, net212741, net212792, net212824,
         net212826, net212840, net212842, net212871, net212874, net212877,
         net212881, net212883, net212886, net212888, net212891, net212893,
         net212900, net212902, net212906, net212909, net212911, net212914,
         net212916, net212920, net212921, net212927, net212928, net212951,
         net212954, net212970, net212971, net212989, net212991, net212999,
         net213000, net213005, net213006, net213012, net213022, net213070,
         net213072, net213111, net213127, net213138, net213140, net213141,
         net213142, net213149, net213152, net213177, net213178, net213229,
         net213244, net213251, net213272, net213275, net213311, net213330,
         net213331, net213332, net213333, net213359, net213364, net213367,
         net213373, net213374, net213375, net213380, net213381, net213383,
         net213410, net213411, net213441, net213473, net213508, net213513,
         net213527, net213528, net213529, net213532, net213533, net213534,
         net213541, net213542, net213543, net213547, net213548, net213553,
         net213555, net213556, net213557, net213560, net213562, net213565,
         net213566, net213567, net213570, net213571, net213572, net213574,
         net213575, net213576, net213577, net213578, net213579, net213581,
         net213592, net213593, net213594, net213598, net213604, net213605,
         net213607, net213608, net213609, net213611, net213612, net213634,
         net213639, net213680, net213683, net213684, net213692, net213701,
         net213702, net213703, net213704, net213705, net213706, net213707,
         net213711, net213712, net213716, net213718, net213722, net213725,
         net213726, net213730, net213732, net213734, net213736, net213737,
         net213738, net213740, net213743, net213745, net213749, net213750,
         net213752, net213753, net213754, net213758, net213759, net213761,
         net213762, net213763, net213764, net213766, net213767, net213769,
         net213770, net213772, net213773, net213775, net213776, net213778,
         net213779, net213780, net213782, net213786, net213787, net213790,
         net213792, net213795, net213797, net213801, net213802, net213805,
         net213806, net213808, net213830, net213837, net213850, net213851,
         net213852, net213864, net213865, net213866, net213867, net213919,
         net213924, net213925, net213926, net213927, net213969, net213981,
         net213983, net213984, net213988, net213989, net213990, net213992,
         net213993, net213994, net213995, net213997, net214019, net214020,
         net214022, net214024, net214025, net214033, net214038, net214039,
         net214057, net214059, net214072, net214073, net214077, net214078,
         net214083, net214084, net214085, net214086, net214087, net214089,
         net214092, net214101, net214103, net214145, net214147, net214152,
         net214172, net214173, net214219, net214224, net214247, net214288,
         net214289, net214293, net214323, net214324, net214325, net214326,
         net214329, net214330, net214331, net214332, net214334, net214338,
         net214339, net214371, net214372, net214376, net214384, net214385,
         net214387, net214391, net214427, net214428, net214429, net214433,
         net214434, net214456, net214457, net214459, net214476, net214477,
         net214478, net214479, net214486, net214487, net214489, net214536,
         net214538, net214549, net214551, net214568, net214571, net214583,
         net214584, net214586, net214588, net214603, net214610, net214611,
         net214612, net214617, net214619, net214620, net214660, net214661,
         net214705, net214710, net214711, net214713, net214716, net214720,
         net214726, net214728, net214730, net214731, net214732, net214747,
         net214758, net214784, net214785, net214792, net214793, net214804,
         net214830, net214834, net214840, net214846, net214853, net214863,
         net214921, net214922, net214926, net214954, net214955, net214963,
         net214964, net214971, net214972, net214974, net214978, net214979,
         net214983, net214984, net215001, net215014, net215022, net215023,
         net215024, net215057, net215058, net215059, net215061, net215062,
         net215064, net215072, net215073, net215089, net215090, net215111,
         net215112, net215114, net215121, net215122, net215124, net215126,
         net215127, net215129, net215175, net215176, net215199, net215204,
         net215206, net215209, net215211, net215212, net215218, net215224,
         net215232, net215245, net215252, net215256, net215275, net215277,
         net215279, net215282, net215287, net215294, net215295, net215296,
         net215298, net215300, net215301, net215307, net215316, net215318,
         net215320, net215324, net215325, net215327, net215328, net215334,
         net215335, net215347, net215357, net215360, net215363, net215414,
         net215416, net215421, net215424, net215431, net215434, net215468,
         net215471, net215475, net215476, net215477, net215478, net215491,
         net215492, net215493, net215494, net215499, net215516, net215517,
         net215518, net215519, net215530, net215565, net215566, net215568,
         net215569, net215571, net215576, net215581, net215582, net215583,
         net215589, net215590, net215591, net215593, net215595, net215635,
         net215636, net215661, net215662, net215663, net215667, net215672,
         net215673, net215674, net215675, net215701, net215709, net215770,
         net215773, net215775, net215776, net215777, net215780, net215781,
         net215782, net215783, net215786, net215790, net215791, net215799,
         net215802, net215805, net215807, net215809, net215812, net215814,
         net215846, net215848, net215853, net215913, net215919, net215920,
         net216001, net216008, net216019, net216020, net216022, net216052,
         net216063, net216064, net216092, net216097, net216117, net216124,
         net216126, net216128, net216129, net216135, net216190, net216191,
         net216192, net216193, net216196, net216198, net216200, net216202,
         net216203, net216211, net216212, net216213, net216217, net216219,
         net216220, net216221, net216222, net216251, net216256, net216259,
         net216277, net216279, net216281, net216283, net216284, net216285,
         net216306, net216327, net216328, net216329, net216330, net216332,
         net216334, net216388, net216392, net216393, net216394, net216400,
         net216436, net216439, net216517, net216520, net216522, net216523,
         net216565, net216566, net216567, net216568, net216569, net216571,
         net216573, net216574, net216575, net216576, net216579, net216584,
         net216587, net216620, net216622, net216627, net216632, net216644,
         net216645, net216649, net216650, net216653, net216692, net216698,
         net216704, net216710, net216711, net216714, net216716, net216759,
         net216760, net216761, net216782, net216783, net216794, net216795,
         net216796, net216811, net216819, net216835, net216839, net216840,
         net216841, net216842, net216843, net216844, net216855, net216856,
         net216885, net216925, net216926, net216927, net216928, net216929,
         net216932, net216934, net216935, net216936, net216941, net216943,
         net216944, net216945, net216947, net216958, net216960, net216965,
         net216968, net216979, net216985, net216987, net216998, net217000,
         net217001, net217027, net217029, net217030, net217031, net217069,
         net217070, net217071, net217072, net217075, net217077, net217082,
         net217083, net217088, net217091, net217092, net217094, net217106,
         net217118, net217121, net217122, net217133, net217141, net217142,
         net217169, net217179, net217182, net217228, net217233, net217235,
         net217236, net217238, net217240, net217242, net217244, net217258,
         net217259, net217260, net217261, net217264, net217267, net217271,
         net217273, net217274, net217275, net217278, net217281, net217282,
         net217283, net217284, net217285, net217287, net217288, net217295,
         net217298, net217299, net217340, net217344, net217346, net217348,
         net217356, net217360, net217361, net217362, net217365, net217376,
         net217395, net217396, net217403, net217408, net217414, net217427,
         net217431, net217433, net217438, net217439, net217442, net217445,
         net217464, net217478, net217497, net217506, net217512, net217517,
         net217524, net217526, net217529, net217541, net217545, net217550,
         net217552, net217557, net217584, net217608, net217621, net217630,
         net217631, net217654, net217677, net217732, net217736, net217759,
         net217761, net217771, net217779, net217780, net217781, net217782,
         net217783, net217786, net217795, net217796, net217806, net217807,
         net217816, net217817, net217818, net217819, net217838, net217849,
         net217858, net217859, net217860, net217876, net217877, net217878,
         net217897, net217933, net217942, net217943, net217944, net217946,
         net217948, net217950, net217960, net217966, net217972, net217973,
         net217977, net217978, net217979, net217982, net217983, net217984,
         net217988, net217989, net217990, net217993, net217994, net217995,
         net218040, net218041, net218042, net218043, net218054, net218058,
         net218059, net218075, net218076, net218079, net218084, net218089,
         net218090, net218091, net218093, net218096, net218097, net218099,
         net218106, net218114, net218115, net218116, net218124, net218132,
         net218133, net218135, net218136, net218137, net218140, net218142,
         net218143, net218144, net218146, net218149, net218156, net218157,
         net218158, net218165, net218166, net218178, net218206, net218207,
         net218208, net218210, net218212, net218214, net218215, net218217,
         net218219, net218220, net218224, net218232, net218236, net218237,
         net218240, net218241, net218244, net218245, net218251, net218256,
         net218257, net218260, net218261, net218262, net218263, net218266,
         net218267, net218269, net218272, net218273, net218276, net218281,
         net218282, net218284, net218285, net218306, net218308, net218321,
         net218322, net218334, net218352, net218353, net218354, net218362,
         net218367, net218370, net218371, net218378, net218392, net218406,
         net218420, net218428, net218442, net218456, net218470, net218486,
         net218484, net218496, net218514, net218530, net218544, net218540,
         net218538, net218536, net218534, net218554, net218550, net218548,
         net218546, net218566, net218562, net218560, net218558, net218556,
         net218576, net218574, net218604, net218600, net218598, net218614,
         net218610, net218608, net218606, net218628, net218626, net218624,
         net218640, net218639, net218655, net218660, net218659, net218809,
         net218808, net219036, net219054, net219055, net219063, net219065,
         net219120, net219116, net219162, net219178, net219328, net219338,
         net219358, net219368, net219468, net219485, net219497, net219557,
         net219556, net219561, net219569, net219611, net219630, net219641,
         net219656, net219657, net219674, net219673, net219679, net219678,
         net219771, net219770, net219859, net219864, net219874, net219931,
         net219934, net219938, net219965, net220022, net220061, net220079,
         net220099, net220153, net220181, net220199, net220293, net220298,
         net220385, net220394, net220396, net220397, net220410, net220496,
         net220521, net214879, net218268, net218238, net218234, net219220,
         net216210, net216207, net216206, net216205, net216096, net216095,
         net215813, net212687, net212404, net218110, net217246, net218235,
         net218233, net218148, net218147, net218145, net217294, net217293,
         net217292, net217291, net215798, net215586, net215585, net215584,
         net215346, net215344, net215342, net212127, net212113, net212099,
         net213756, net213755, net213751, net213443, net213442, net213439,
         net213201, net223182, net223234, net223412, net223422, net223484,
         net223505, net223581, net223586, net223617, net223689, net223706,
         net223819, net223932, net224032, net224078, net223271, net223270,
         net219978, net215792, net215784, net215343, net215337, net214877,
         net218100, net213409, net213234, net213232, net216282, net212641,
         net213239, net213238, net219526, net216978, net216767, net216763,
         net216585, net216226, net214969, net214968, net214864, net214961,
         net214960, net214959, net218221, net218174, net218173, net218098,
         net218095, net218094, net217262, net223908, net215308, net214832,
         net214831, net214569, net218105, net218101, net217290, net217109,
         net214727, net214724, net214723, net215322, net215219, net214857,
         net214856, net212452, net214818, net214817, net214721, net219847,
         net216836, net216660, net216578, net216577, net218139, net218057,
         net217230, net217229, net213401, net213400, net213407, net213406,
         net213405, net213404, net213237, net214786, net214546, net214545,
         net214542, net216651, net216647, net219339, net219238, net219237,
         net219236, net216762, net216658, net216657, net216583, net216582,
         net216572, net219746, net212644, net212642, net212640, net215082,
         net215081, net215078, net215076, net215075, net215447, net215446,
         net215445, net215216, net215215, net215214, net214967, net213700,
         net220149, net215339, net215210, net216776, net216775, net216774,
         net216773, net217863, net213729, net213724, net213719, net213589,
         net213587, net213586, net213233, net219976, net217086, net217085,
         net217084, net217081, net216652, net218271, net218239, net218216,
         net220033, net218270, net216094, net215797, net223718, net215338,
         net215336, net215332, net215331, net215330, net215329, net215217,
         net219540, net219539, net214174, net213982, net213892, net213891,
         net213889, net213888, net213887, net213588, net212650, net215354,
         net215351, net215350, net219749, net212733, net223531, net220019,
         net218109, net218065, net218063, net218061, net218060, net217237,
         net217231, net219781, net216209, net216208, net216018, net215796,
         net215793, net215668, net219713, net219494, net219256, net217232,
         net217079, net217078, net216834, net216833, net216832, net216831,
         net216830, net216777, net216771, net216770, net216769, net216768,
         net216648, net216646, net214541, net214539, net214179, net214178,
         net214175, net215102, net215100, net215099, net223874, net215310,
         net215088, net215087, net215085, net215084, net215083, net214973,
         net214570, net223712, net215096, net215094, net219336, net216017,
         net216016, net215811, net215810, net215808, net215806, net215669,
         net217790, net219530, net219429, net214815, net214814, net214812,
         net214811, net214810, net214717, net214715, net214461, net219069,
         net214809, net214808, net214797, net214796, net214795, net214794,
         net214543, net214460, net220004, net215213, net215107, net215106,
         net215105, net215104, net215103, net214966, net214855, net213402,
         net213399, net213248, net213242, net218175, net218172, net218171,
         net218170, net218153, net218152, net218151, net218150, net218072,
         net218071, net218070, net218069, net218068, net218067, net218066,
         net217243, net216946, net220046, net213595, net213398, net213397,
         net213394, net223508, net215095, net215093, net215092, net215091,
         net214975, net214714, net215352, net215349, net215348, net215123,
         net214878, net215101, net215098, net215097, net214970, net214587,
         net218112, net218111, net218104, net218103, net217107, net220449,
         net213606, net213603, net213396, net213395, net213393, net213388,
         net213033, net213031, net213023, net212942, net215302, net215077,
         net215074, net214820, net214819, net214719, net214718, net220395,
         net218339, net218337, net218297, net218277, net217879, net217857,
         net223455, net215666, net215665, net215664, net215587, net215430,
         net215429, net215428, net215427, net215426, net215425, net215353,
         net214958, net241090, net241077, net241076, net241055, net241366,
         net241365, net241364, net241372, net241371, net213522, net213512,
         net213791, net213539, net213538, net213537, net220211, net220210,
         net213408, net213231, net213230, net212925, net213546, net213191,
         net213190, net213804, net213139, net213132, net213131, net213130,
         net213222, net213183, net213472, net213167, net213115, net213438,
         net213437, net213436, net213208, net213207, net213392, net213391,
         net213389, net213384, net213024, net213021, net213019, net213403,
         net213236, net213235, net212930, net241088, net241082, net241074,
         net241071, net212454, net213217, net214093, net214090, net213822,
         net213821, net212419, net212715, net220036, net213818, net213514,
         net213520, net217899, net213551, net213196, net213195, net214924,
         net214668, net215418, net215183, net223123, net223105, net212399,
         net212112, net212111, net212110, net212103, net213583, net213580,
         net213413, net213225, net213041, net213040, net212429, net212428,
         net212418, net220017, net213713, net213597, net213602, net213464,
         net213463, net213181, net218502, net213446, net214389, net214100,
         net216624, net216446, net218480, net212683, net212402, net212401,
         net213469, net213468, net216253, net216072, net213454, net213452,
         net213451, net213193, net213192, net213524, net213523, net213418,
         net213417, net213416, net213415, net213227, net213220, net219068,
         net212648, net212441, net213460, net213458, net213457, net213188,
         net213187, net214394, net214929, net213483, net213481, net213113,
         net213488, net213486, net213165, net213495, net213493, net213491,
         net213129, net213386, net213382, net213250, net213249, net212948,
         net212947, net212944, net212732, net213870, net213448, net213197,
         net213596, net213247, net213246, net213245, net213243, net213241,
         net213240, net213036, net212935, net216623, net216444, net216441,
         net213833, net223121, net223119, net223089, net223090, net219445,
         net218476, net212398, net212397, net212389, net212945, net212724,
         net212723, net212722, net212721, net212720, net212719, net212647,
         net217136, net217280, net217183, net217140, net217131, net217130,
         net217127, net217124, net223812, net218552, net213832, net213826,
         net213824, net213823, net213516, net213515, net213511, net220146,
         net220145, net213020, net213018, net213016, net213015, net213014,
         net213013, net212946, net211944, net214928, net214666, net214665,
         net214663, net214662, net214395, net215417, net215181, net215180,
         net215178, net215177, net214930, net217970, net217028, net215855,
         net215850, net215644, net213465, net213462, net213461, net213189,
         net213186, net213185, net213484, net213482, net213173, net213171,
         net213489, net213487, net213485, net213116, net213114, net213112,
         net213494, net213492, net213490, net213168, net213166, net213164,
         net218542, net213816, net213814, net213521, net213519, net213470,
         net213467, net213466, net213184, net213182, net213180, net213453,
         net213450, net213449, net213198, net212795, net212794, net213211,
         net223498, net223481, net223126, net223125, net223124, net223109,
         net223104, net223100, net223098, net223009, net212405, net212403,
         net212105, net220060, net215854, net215849, net215643, net215642,
         net215641, net215640, net215423, net215422, net215186, net215185,
         net215184, net213042, net213039, net213038, net212936, net212934,
         net212932, net223607, net223606, net223578, net223577, net218658,
         net212104, net212100, net212097, net213414, net213226, net213054,
         net213050, net212919, net212918, net213046, net213045, net212923,
         net213422, net213421, net213215, net224038, net213447, net213445,
         net213444, net213206, net213203, net218414, net216962, net216800,
         net216252, net216070, net216069, net216068, net216067, net215856,
         net214393, net214098, net214097, net214096, net214095, net213834,
         net219990, net218400, net213435, net213434, net213433, net213431,
         net213430, net213213, net213205, net213204, net213202, net223487,
         net213429, net213426, net213212, net213209, net218164, net218578,
         net218434, net218161, net218568, net218160, net218159, net218083,
         net218082, net218081, net217276, net217139, net217138, net217135,
         net213813, net213812, net213810, net213809, net213518, net213517,
         net220011, net219412, net212432, net212431, net212430, net212423,
         net212416, net212415, net212414, net212413, net212390, net212122,
         net219974, net213480, net213479, net213478, net213477, net213475,
         net213176, net213174, net213172, net213170, net213169, net213035,
         net213034, net213459, net213456, net213455, net213194, net212899,
         net212713, net224071, net213428, net213427, net213424, net213218,
         net213216, net213214, net213210, net213047, net213044, net213043,
         net212931, net212929, net220068, net213053, net213052, net213049,
         net213048, net212926, net212924, net212922, net216443, net216442,
         net216258, net216257, net216075, net216074, net216073, net216961,
         net216799, net216798, net216797, net216631, net216630, net216628,
         net216449, net216448, net216447, net217126, net217125, net216967,
         net216966, net216803, net216802, net216801, net224024, net219464,
         net219463, net219422, net219421, net219357, net219333, net212718,
         net212717, net212714, net212711, net212710, net212709, net212708,
         net212707, net212445, net212440, net212439, net212424, net212422,
         net219933, net219693, net219504, net219503, net213600, net213030,
         net213029, net213028, net213027, net213026, net213025, net213017,
         net212941, net212940, net212939, net212938, net212933, net212731,
         net212643, net213423, net213420, net213419, net213223, net213221,
         net213219, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894;

  INV_X4 U3179 ( .A(n3158), .ZN(n509) );
  DLH_X2 sel_reg ( .G(n3990), .D(n509), .Q(sel) );
  NOR2_X2 U3195 ( .A1(net218109), .A2(net217242), .ZN(n3657) );
  NAND2_X2 U3196 ( .A1(b[1]), .A2(a[2]), .ZN(n3596) );
  INV_X16 U3197 ( .A(net218558), .ZN(n3301) );
  INV_X1 U3198 ( .A(net213246), .ZN(n3194) );
  NAND2_X4 U3199 ( .A1(n7324), .A2(n7325), .ZN(n7395) );
  OAI21_X4 U3200 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6732) );
  NAND2_X4 U3201 ( .A1(n6510), .A2(n6715), .ZN(n6378) );
  NAND2_X4 U3202 ( .A1(n4834), .A2(n4835), .ZN(n4755) );
  NAND2_X4 U3203 ( .A1(n4142), .A2(n4141), .ZN(n4150) );
  INV_X1 U3204 ( .A(n6320), .ZN(n6324) );
  INV_X8 U3205 ( .A(n6168), .ZN(n6054) );
  INV_X1 U3206 ( .A(net216067), .ZN(net219556) );
  INV_X4 U3207 ( .A(n5082), .ZN(n5007) );
  INV_X4 U3208 ( .A(net215075), .ZN(net215077) );
  NAND2_X4 U3209 ( .A1(n3889), .A2(n5548), .ZN(n5626) );
  NAND2_X4 U3210 ( .A1(n5725), .A2(n5724), .ZN(n5766) );
  NAND2_X4 U3211 ( .A1(net218042), .A2(net218043), .ZN(net218040) );
  INV_X2 U3212 ( .A(n5862), .ZN(n5859) );
  INV_X4 U3213 ( .A(net215793), .ZN(net220521) );
  INV_X4 U3214 ( .A(net216762), .ZN(net219339) );
  NAND2_X2 U3215 ( .A1(net213553), .A2(net213556), .ZN(net214330) );
  NAND2_X2 U3216 ( .A1(n6012), .A2(n5972), .ZN(n3166) );
  INV_X2 U3217 ( .A(n5623), .ZN(n5553) );
  INV_X8 U3218 ( .A(net215668), .ZN(net215665) );
  NAND2_X4 U3219 ( .A1(n6723), .A2(n6722), .ZN(n6767) );
  XNOR2_X2 U3220 ( .A(n5939), .B(n5800), .ZN(n3966) );
  INV_X2 U3221 ( .A(n5939), .ZN(n5801) );
  OAI21_X1 U3222 ( .B1(n5805), .B2(n3786), .A(n3572), .ZN(n5675) );
  CLKBUF_X3 U3223 ( .A(n5956), .Z(n3931) );
  NAND2_X4 U3224 ( .A1(n6679), .A2(n6678), .ZN(n6940) );
  INV_X8 U3225 ( .A(net212951), .ZN(n3524) );
  NAND2_X2 U3226 ( .A1(n5522), .A2(n5521), .ZN(n5278) );
  NAND2_X2 U3227 ( .A1(net216022), .A2(net216019), .ZN(n5266) );
  INV_X2 U3228 ( .A(n7396), .ZN(n7397) );
  NAND2_X2 U3229 ( .A1(n3978), .A2(n5298), .ZN(n5425) );
  INV_X2 U3230 ( .A(n5713), .ZN(n5711) );
  NAND2_X4 U3231 ( .A1(n7300), .A2(n7299), .ZN(n7147) );
  NAND2_X4 U3232 ( .A1(n6534), .A2(n6532), .ZN(n6350) );
  INV_X4 U3233 ( .A(net213555), .ZN(n3511) );
  INV_X4 U3234 ( .A(n6236), .ZN(n6237) );
  INV_X8 U3235 ( .A(n5285), .ZN(n5541) );
  INV_X4 U3236 ( .A(n7512), .ZN(n7342) );
  INV_X2 U3237 ( .A(net213751), .ZN(net213754) );
  INV_X2 U3238 ( .A(net213775), .ZN(n3559) );
  INV_X8 U3239 ( .A(n3864), .ZN(net214428) );
  INV_X2 U3240 ( .A(n7516), .ZN(n7520) );
  INV_X2 U3241 ( .A(n3933), .ZN(n7315) );
  XNOR2_X1 U3242 ( .A(net212842), .B(n3767), .ZN(n3938) );
  NAND2_X4 U3243 ( .A1(n6552), .A2(n6551), .ZN(n6738) );
  INV_X8 U3244 ( .A(n3732), .ZN(n3731) );
  NAND2_X4 U3245 ( .A1(n3219), .A2(n3220), .ZN(n3222) );
  INV_X8 U3246 ( .A(net213212), .ZN(net213210) );
  OAI21_X4 U3247 ( .B1(n3317), .B2(n6048), .A(n6167), .ZN(n6168) );
  OAI21_X4 U3248 ( .B1(net213231), .B2(net213230), .A(net220211), .ZN(n3161)
         );
  INV_X2 U3249 ( .A(n5345), .ZN(n3162) );
  CLKBUF_X3 U3250 ( .A(net216200), .Z(n3163) );
  NAND2_X2 U3251 ( .A1(n3164), .A2(n3165), .ZN(n3167) );
  NAND2_X2 U3252 ( .A1(n3166), .A2(n3167), .ZN(n5857) );
  INV_X4 U3253 ( .A(n6012), .ZN(n3164) );
  INV_X2 U3254 ( .A(n5972), .ZN(n3165) );
  NAND2_X2 U3255 ( .A1(n5722), .A2(n3169), .ZN(n3170) );
  NAND2_X2 U3256 ( .A1(n3168), .A2(n5721), .ZN(n3171) );
  NAND2_X2 U3257 ( .A1(n3170), .A2(n3171), .ZN(n3975) );
  INV_X1 U3258 ( .A(n5722), .ZN(n3168) );
  INV_X4 U3259 ( .A(n5721), .ZN(n3169) );
  INV_X4 U3260 ( .A(n5707), .ZN(n3172) );
  NAND2_X4 U3261 ( .A1(b[17]), .A2(a[2]), .ZN(n5972) );
  INV_X8 U3262 ( .A(n3693), .ZN(n3689) );
  INV_X4 U3263 ( .A(net216205), .ZN(net216096) );
  NAND2_X4 U3264 ( .A1(net216001), .A2(net215790), .ZN(n5398) );
  INV_X4 U3265 ( .A(net213593), .ZN(n3748) );
  NAND2_X2 U3266 ( .A1(n6712), .A2(n6710), .ZN(n6386) );
  INV_X4 U3267 ( .A(net214588), .ZN(net214583) );
  INV_X4 U3268 ( .A(n5814), .ZN(n5812) );
  INV_X2 U3269 ( .A(net215431), .ZN(n3608) );
  NAND2_X1 U3270 ( .A1(n5356), .A2(n3806), .ZN(n3173) );
  NAND2_X4 U3271 ( .A1(n3294), .A2(n3295), .ZN(net213732) );
  NAND2_X2 U3272 ( .A1(net213734), .A2(net213574), .ZN(n3294) );
  NAND2_X4 U3273 ( .A1(net215666), .A2(net215584), .ZN(net223271) );
  NAND2_X4 U3274 ( .A1(net213436), .A2(net213437), .ZN(net213207) );
  NAND2_X4 U3275 ( .A1(n3780), .A2(n5798), .ZN(n5669) );
  NAND2_X4 U3276 ( .A1(net212795), .A2(net212794), .ZN(net212634) );
  NAND2_X2 U3277 ( .A1(n6496), .A2(n6495), .ZN(n6700) );
  NAND2_X4 U3278 ( .A1(net216576), .A2(n3693), .ZN(net216760) );
  INV_X2 U3279 ( .A(net216576), .ZN(net216575) );
  NAND2_X2 U3280 ( .A1(net218054), .A2(net217295), .ZN(n3585) );
  AOI21_X4 U3281 ( .B1(n6696), .B2(n6697), .A(n3878), .ZN(n6886) );
  AOI21_X4 U3282 ( .B1(net216573), .B2(net216574), .A(net216575), .ZN(n5123)
         );
  NAND2_X2 U3283 ( .A1(net216226), .A2(n3675), .ZN(net216763) );
  INV_X16 U3284 ( .A(b[1]), .ZN(n3298) );
  INV_X2 U3285 ( .A(n5294), .ZN(n3970) );
  INV_X2 U3286 ( .A(net212925), .ZN(net212923) );
  NAND2_X4 U3287 ( .A1(net214456), .A2(net214457), .ZN(n6418) );
  INV_X2 U3288 ( .A(n6710), .ZN(n6711) );
  NAND2_X4 U3289 ( .A1(n3813), .A2(n3814), .ZN(n3815) );
  INV_X1 U3290 ( .A(n6427), .ZN(n6431) );
  CLKBUF_X2 U3291 ( .A(net218104), .Z(n3174) );
  NAND2_X4 U3292 ( .A1(n6369), .A2(n6370), .ZN(n6512) );
  NAND2_X2 U3293 ( .A1(n6520), .A2(n6519), .ZN(n6362) );
  NAND2_X4 U3294 ( .A1(net214832), .A2(net214569), .ZN(n3688) );
  XNOR2_X2 U3295 ( .A(n5965), .B(net215316), .ZN(n3883) );
  NAND2_X4 U3296 ( .A1(net215217), .A2(net214969), .ZN(net215328) );
  INV_X4 U3297 ( .A(net213566), .ZN(n3448) );
  INV_X4 U3298 ( .A(net213213), .ZN(net213209) );
  NAND2_X4 U3299 ( .A1(n6512), .A2(n6720), .ZN(n6373) );
  NAND2_X2 U3300 ( .A1(n6515), .A2(n6514), .ZN(n6368) );
  NAND2_X4 U3301 ( .A1(net212951), .A2(net212655), .ZN(n7108) );
  INV_X2 U3302 ( .A(net216209), .ZN(net216568) );
  BUF_X8 U3303 ( .A(net216587), .Z(net219497) );
  INV_X2 U3304 ( .A(n3687), .ZN(n3257) );
  NAND2_X4 U3305 ( .A1(net215185), .A2(net215186), .ZN(net215184) );
  NAND2_X4 U3306 ( .A1(n7157), .A2(n7158), .ZN(n7253) );
  OAI21_X4 U3307 ( .B1(n4163), .B2(n4737), .A(n4736), .ZN(n4156) );
  NAND2_X1 U3308 ( .A1(n3315), .A2(n5385), .ZN(n3175) );
  NAND2_X1 U3309 ( .A1(net212933), .A2(net213038), .ZN(n3178) );
  NAND2_X2 U3310 ( .A1(n3176), .A2(n3177), .ZN(n3179) );
  NAND2_X2 U3311 ( .A1(n3178), .A2(n3179), .ZN(net219693) );
  INV_X4 U3312 ( .A(net212933), .ZN(n3176) );
  INV_X2 U3313 ( .A(net213038), .ZN(n3177) );
  NOR2_X4 U3314 ( .A1(n3180), .A2(n3181), .ZN(n3182) );
  NOR2_X4 U3315 ( .A1(n3182), .A2(net213226), .ZN(net212919) );
  INV_X4 U3316 ( .A(net213413), .ZN(n3180) );
  INV_X2 U3317 ( .A(net213225), .ZN(n3181) );
  NAND2_X2 U3318 ( .A1(net213454), .A2(net213455), .ZN(n3185) );
  NAND2_X4 U3319 ( .A1(n3183), .A2(n3184), .ZN(n3186) );
  NAND2_X4 U3320 ( .A1(n3185), .A2(n3186), .ZN(net213451) );
  INV_X4 U3321 ( .A(net213454), .ZN(n3183) );
  INV_X4 U3322 ( .A(net213455), .ZN(n3184) );
  NAND2_X2 U3323 ( .A1(net213419), .A2(net213222), .ZN(n3189) );
  NAND2_X4 U3324 ( .A1(n3187), .A2(n3188), .ZN(n3190) );
  NAND2_X4 U3325 ( .A1(n3189), .A2(n3190), .ZN(net213417) );
  INV_X4 U3326 ( .A(net213419), .ZN(n3187) );
  INV_X2 U3327 ( .A(net213222), .ZN(n3188) );
  NAND2_X2 U3328 ( .A1(n3315), .A2(n5385), .ZN(n3210) );
  INV_X2 U3329 ( .A(net213227), .ZN(net213226) );
  NAND2_X4 U3330 ( .A1(net213450), .A2(net213451), .ZN(net212794) );
  INV_X2 U3331 ( .A(net213417), .ZN(net213415) );
  INV_X2 U3332 ( .A(net212940), .ZN(net212939) );
  INV_X1 U3333 ( .A(net219539), .ZN(net214173) );
  OAI21_X1 U3334 ( .B1(n5726), .B2(n5761), .A(n5762), .ZN(n5727) );
  NAND2_X1 U3335 ( .A1(n5764), .A2(n5762), .ZN(n5589) );
  XNOR2_X2 U3336 ( .A(net213438), .B(net213439), .ZN(net213437) );
  INV_X4 U3337 ( .A(net213208), .ZN(net213204) );
  INV_X1 U3338 ( .A(n6514), .ZN(n6518) );
  INV_X2 U3339 ( .A(n6519), .ZN(n6523) );
  NAND2_X4 U3340 ( .A1(n6322), .A2(n6519), .ZN(n6198) );
  OAI21_X1 U3341 ( .B1(net212696), .B2(n3363), .A(net212429), .ZN(net212991)
         );
  OAI21_X2 U3342 ( .B1(net212696), .B2(n3363), .A(net212697), .ZN(net212428)
         );
  NAND2_X4 U3343 ( .A1(n6968), .A2(n6967), .ZN(net213375) );
  NAND2_X2 U3344 ( .A1(n6623), .A2(n6624), .ZN(n6833) );
  NAND2_X1 U3345 ( .A1(n5685), .A2(n5684), .ZN(n3571) );
  INV_X1 U3346 ( .A(n7241), .ZN(n7243) );
  INV_X2 U3347 ( .A(n6895), .ZN(n6899) );
  INV_X4 U3348 ( .A(net212929), .ZN(net219673) );
  NAND2_X4 U3349 ( .A1(net213020), .A2(n3243), .ZN(net213018) );
  OAI21_X2 U3350 ( .B1(n4748), .B2(n4824), .A(n4825), .ZN(n4749) );
  NOR2_X1 U3351 ( .A1(net220396), .A2(n3620), .ZN(net218339) );
  OAI21_X4 U3352 ( .B1(net212732), .B2(net212733), .A(net219749), .ZN(
        net212642) );
  INV_X2 U3353 ( .A(net216572), .ZN(net216571) );
  INV_X1 U3354 ( .A(n5222), .ZN(n5227) );
  NAND2_X4 U3355 ( .A1(net214818), .A2(net214719), .ZN(net215073) );
  NAND2_X4 U3356 ( .A1(net215075), .A2(net215074), .ZN(net214719) );
  NAND2_X4 U3357 ( .A1(net216660), .A2(net216926), .ZN(net216925) );
  XNOR2_X2 U3358 ( .A(n4717), .B(n4986), .ZN(n4718) );
  NAND2_X4 U3359 ( .A1(n7248), .A2(net212902), .ZN(n7501) );
  NAND2_X4 U3360 ( .A1(n5505), .A2(n5779), .ZN(n5651) );
  INV_X4 U3361 ( .A(n6968), .ZN(n6965) );
  XNOR2_X2 U3362 ( .A(n7025), .B(net212653), .ZN(n3766) );
  INV_X2 U3363 ( .A(n3530), .ZN(n3191) );
  INV_X4 U3364 ( .A(n7100), .ZN(n7044) );
  AOI21_X2 U3365 ( .B1(b[27]), .B2(n7032), .A(n3389), .ZN(n7066) );
  NAND2_X4 U3366 ( .A1(n7013), .A2(n7012), .ZN(n6963) );
  NAND2_X4 U3367 ( .A1(net212428), .A2(net212429), .ZN(net212694) );
  OAI21_X2 U3368 ( .B1(n3530), .B2(n3531), .A(net212703), .ZN(n3529) );
  NAND2_X2 U3369 ( .A1(n6803), .A2(n6804), .ZN(n3192) );
  NAND2_X2 U3370 ( .A1(n6790), .A2(n6791), .ZN(n3193) );
  NAND2_X2 U3371 ( .A1(n6618), .A2(n6617), .ZN(n3195) );
  NAND2_X2 U3372 ( .A1(n6618), .A2(n6617), .ZN(n6955) );
  NAND2_X2 U3373 ( .A1(n5935), .A2(n3310), .ZN(n6050) );
  XNOR2_X2 U3374 ( .A(n3655), .B(net218065), .ZN(n3196) );
  XNOR2_X2 U3375 ( .A(n5973), .B(n3777), .ZN(n5974) );
  NAND2_X4 U3376 ( .A1(n5975), .A2(n5974), .ZN(net214731) );
  CLKBUF_X2 U3377 ( .A(n5649), .Z(n3197) );
  INV_X2 U3378 ( .A(net213242), .ZN(n3198) );
  INV_X4 U3379 ( .A(n3198), .ZN(n3199) );
  OAI21_X4 U3380 ( .B1(n3508), .B2(n3509), .A(net213551), .ZN(net213195) );
  INV_X4 U3381 ( .A(net213764), .ZN(n3508) );
  INV_X2 U3382 ( .A(net213196), .ZN(net213192) );
  XNOR2_X2 U3383 ( .A(n7336), .B(n7335), .ZN(n3200) );
  OAI21_X4 U3384 ( .B1(n3890), .B2(n7105), .A(n7104), .ZN(n7111) );
  NAND2_X4 U3385 ( .A1(n6254), .A2(n6253), .ZN(n6427) );
  INV_X2 U3386 ( .A(n6414), .ZN(n6416) );
  INV_X2 U3387 ( .A(n5259), .ZN(n5256) );
  XNOR2_X2 U3388 ( .A(n6797), .B(n6893), .ZN(n3201) );
  INV_X4 U3389 ( .A(n6893), .ZN(n6798) );
  INV_X2 U3390 ( .A(net215127), .ZN(n3868) );
  NAND2_X4 U3391 ( .A1(net215791), .A2(net215790), .ZN(n5688) );
  NOR3_X4 U3392 ( .A1(net212660), .A2(n7391), .A3(n7390), .ZN(n7392) );
  INV_X4 U3393 ( .A(n4918), .ZN(n3202) );
  NAND2_X2 U3394 ( .A1(net215214), .A2(net215215), .ZN(net215327) );
  NAND2_X2 U3395 ( .A1(net215475), .A2(net215476), .ZN(n5580) );
  NAND2_X1 U3396 ( .A1(n5581), .A2(net215476), .ZN(n5444) );
  XNOR2_X2 U3397 ( .A(n6563), .B(n6562), .ZN(n3203) );
  NAND2_X4 U3398 ( .A1(n6728), .A2(n6731), .ZN(n6562) );
  XNOR2_X2 U3399 ( .A(n5669), .B(n5668), .ZN(n3204) );
  AND2_X2 U3400 ( .A1(n7050), .A2(n6451), .ZN(n3205) );
  AND2_X4 U3401 ( .A1(net218094), .A2(net218098), .ZN(n3206) );
  INV_X8 U3402 ( .A(net217109), .ZN(net218072) );
  NAND2_X4 U3403 ( .A1(n6542), .A2(n6541), .ZN(n6344) );
  NAND2_X4 U3404 ( .A1(n5784), .A2(n5783), .ZN(n5658) );
  NAND2_X4 U3405 ( .A1(n4055), .A2(n4054), .ZN(net218257) );
  NAND2_X4 U3406 ( .A1(net217246), .A2(net217732), .ZN(n3288) );
  AOI21_X4 U3407 ( .B1(n5361), .B2(n5246), .A(n5245), .ZN(n5247) );
  NAND2_X4 U3408 ( .A1(n5355), .A2(n5115), .ZN(n5224) );
  INV_X8 U3409 ( .A(n4151), .ZN(n4137) );
  NAND2_X4 U3410 ( .A1(n4793), .A2(n4792), .ZN(n4731) );
  NAND2_X4 U3411 ( .A1(net216219), .A2(net216393), .ZN(n3654) );
  OAI21_X4 U3412 ( .B1(n3321), .B2(n3973), .A(n5956), .ZN(n5957) );
  INV_X2 U3413 ( .A(net216210), .ZN(net216095) );
  NAND2_X4 U3414 ( .A1(net215813), .A2(net216020), .ZN(net216210) );
  NAND2_X4 U3415 ( .A1(n4883), .A2(net216932), .ZN(n3746) );
  NAND2_X4 U3416 ( .A1(n4886), .A2(n4885), .ZN(n4883) );
  INV_X8 U3417 ( .A(net215796), .ZN(n3603) );
  NAND2_X4 U3418 ( .A1(n5961), .A2(net215363), .ZN(n5817) );
  NAND2_X4 U3419 ( .A1(n6721), .A2(n6720), .ZN(n6723) );
  INV_X8 U3420 ( .A(n5912), .ZN(n3764) );
  NAND2_X4 U3421 ( .A1(n5616), .A2(n5618), .ZN(n5429) );
  NAND2_X4 U3422 ( .A1(n5822), .A2(n5913), .ZN(net215775) );
  INV_X4 U3423 ( .A(net213557), .ZN(n3219) );
  NAND2_X4 U3424 ( .A1(n6782), .A2(n6783), .ZN(net213441) );
  AND2_X2 U3425 ( .A1(n3482), .A2(net213441), .ZN(n3207) );
  NAND2_X4 U3426 ( .A1(net213753), .A2(net213754), .ZN(net213750) );
  NAND2_X4 U3427 ( .A1(net223874), .A2(net215085), .ZN(n3639) );
  NAND2_X4 U3428 ( .A1(n6671), .A2(n6670), .ZN(n6873) );
  AND2_X4 U3429 ( .A1(n3431), .A2(net213600), .ZN(n3208) );
  NAND2_X4 U3430 ( .A1(net212947), .A2(net212948), .ZN(n3476) );
  NAND2_X4 U3431 ( .A1(net212938), .A2(net212940), .ZN(net213029) );
  AOI21_X4 U3432 ( .B1(net212938), .B2(net213030), .A(net212939), .ZN(
        net220079) );
  NAND2_X4 U3433 ( .A1(net212645), .A2(net212641), .ZN(n3540) );
  INV_X8 U3434 ( .A(net215576), .ZN(net215571) );
  NAND2_X4 U3435 ( .A1(net215434), .A2(net215335), .ZN(net215576) );
  INV_X4 U3436 ( .A(n5354), .ZN(n5358) );
  NAND2_X4 U3437 ( .A1(net213442), .A2(net213201), .ZN(net213756) );
  NAND2_X1 U3438 ( .A1(n5622), .A2(n5624), .ZN(n5554) );
  NAND2_X2 U3439 ( .A1(n5470), .A2(n5473), .ZN(n5346) );
  NAND2_X4 U3440 ( .A1(net217294), .A2(net218106), .ZN(net218208) );
  INV_X2 U3441 ( .A(n7130), .ZN(n7128) );
  NAND2_X1 U3442 ( .A1(n3615), .A2(net218276), .ZN(n3209) );
  NAND2_X4 U3443 ( .A1(net213780), .A2(n6929), .ZN(net213543) );
  NAND2_X4 U3444 ( .A1(n5660), .A2(n5659), .ZN(n5662) );
  INV_X2 U3445 ( .A(n6307), .ZN(n3953) );
  NAND2_X2 U3446 ( .A1(n6164), .A2(n6325), .ZN(n6059) );
  NAND2_X4 U3447 ( .A1(net217291), .A2(net217292), .ZN(net217288) );
  NAND2_X2 U3448 ( .A1(n6026), .A2(n5962), .ZN(n5816) );
  INV_X8 U3449 ( .A(n5962), .ZN(n6022) );
  INV_X2 U3450 ( .A(net218135), .ZN(net218139) );
  NAND2_X4 U3451 ( .A1(net218151), .A2(n3569), .ZN(net217107) );
  NAND2_X2 U3452 ( .A1(n3850), .A2(net214339), .ZN(n3843) );
  OAI21_X4 U3453 ( .B1(n6498), .B2(n6497), .A(n6705), .ZN(n6577) );
  NAND2_X2 U3454 ( .A1(net214152), .A2(net214147), .ZN(n6576) );
  NAND2_X4 U3455 ( .A1(n7238), .A2(n7239), .ZN(n7186) );
  NAND2_X4 U3456 ( .A1(n4041), .A2(net220153), .ZN(n4043) );
  OAI21_X2 U3457 ( .B1(net241090), .B2(net241055), .A(net212641), .ZN(
        net212146) );
  INV_X1 U3458 ( .A(n5920), .ZN(n5924) );
  INV_X4 U3459 ( .A(net215784), .ZN(net219978) );
  INV_X2 U3460 ( .A(n6793), .ZN(n3290) );
  NAND2_X2 U3461 ( .A1(net214551), .A2(net214459), .ZN(n3640) );
  INV_X4 U3462 ( .A(n6407), .ZN(n6405) );
  XNOR2_X1 U3463 ( .A(n3731), .B(net215360), .ZN(n3729) );
  INV_X2 U3464 ( .A(n4054), .ZN(n4037) );
  INV_X8 U3465 ( .A(n4963), .ZN(n4970) );
  NAND2_X2 U3466 ( .A1(n6900), .A2(n6901), .ZN(n6772) );
  OAI21_X4 U3467 ( .B1(n3865), .B2(net215122), .A(n3866), .ZN(n3864) );
  NAND2_X2 U3468 ( .A1(n3632), .A2(net214804), .ZN(n3630) );
  INV_X4 U3469 ( .A(net213596), .ZN(net213245) );
  INV_X8 U3470 ( .A(n7413), .ZN(n7303) );
  NAND2_X4 U3471 ( .A1(n7403), .A2(n7401), .ZN(n7317) );
  INV_X4 U3472 ( .A(n6826), .ZN(n6827) );
  NAND2_X1 U3473 ( .A1(net223125), .A2(net223124), .ZN(n3213) );
  NAND2_X4 U3474 ( .A1(n3211), .A2(n3212), .ZN(n3214) );
  NAND2_X2 U3475 ( .A1(n3213), .A2(n3214), .ZN(net223104) );
  INV_X4 U3476 ( .A(net223125), .ZN(n3211) );
  INV_X4 U3477 ( .A(net223124), .ZN(n3212) );
  NAND2_X1 U3478 ( .A1(net213439), .A2(net213443), .ZN(n3217) );
  NAND2_X2 U3479 ( .A1(n3215), .A2(n3216), .ZN(n3218) );
  NAND2_X2 U3480 ( .A1(n3217), .A2(n3218), .ZN(net213755) );
  INV_X4 U3481 ( .A(net213439), .ZN(n3215) );
  INV_X1 U3482 ( .A(net213443), .ZN(n3216) );
  NAND2_X1 U3483 ( .A1(net213557), .A2(net214022), .ZN(n3221) );
  NAND2_X2 U3484 ( .A1(n3221), .A2(n3222), .ZN(net214329) );
  INV_X1 U3485 ( .A(net214022), .ZN(n3220) );
  NAND2_X1 U3486 ( .A1(net215348), .A2(net215210), .ZN(n3225) );
  NAND2_X2 U3487 ( .A1(n3223), .A2(n3224), .ZN(n3226) );
  NAND2_X2 U3488 ( .A1(n3225), .A2(n3226), .ZN(net215339) );
  INV_X4 U3489 ( .A(net215348), .ZN(n3223) );
  INV_X1 U3490 ( .A(net215210), .ZN(n3224) );
  NAND2_X1 U3491 ( .A1(net213391), .A2(net213392), .ZN(n3229) );
  NAND2_X2 U3492 ( .A1(n3227), .A2(n3228), .ZN(n3230) );
  NAND2_X2 U3493 ( .A1(n3229), .A2(n3230), .ZN(n3541) );
  INV_X4 U3494 ( .A(net213391), .ZN(n3227) );
  INV_X4 U3495 ( .A(net213392), .ZN(n3228) );
  NAND2_X1 U3496 ( .A1(net216016), .A2(net216017), .ZN(n3233) );
  NAND2_X2 U3497 ( .A1(n3231), .A2(n3232), .ZN(n3234) );
  NAND2_X4 U3498 ( .A1(n3233), .A2(n3234), .ZN(n3637) );
  INV_X4 U3499 ( .A(net216016), .ZN(n3231) );
  INV_X2 U3500 ( .A(net216017), .ZN(n3232) );
  NAND2_X2 U3501 ( .A1(n4807), .A2(n4806), .ZN(n3237) );
  NAND2_X4 U3502 ( .A1(n3235), .A2(n3236), .ZN(n3238) );
  NAND2_X4 U3503 ( .A1(n3237), .A2(n3238), .ZN(n4811) );
  INV_X4 U3504 ( .A(n4807), .ZN(n3235) );
  INV_X8 U3505 ( .A(n4806), .ZN(n3236) );
  INV_X8 U3506 ( .A(net223009), .ZN(net223124) );
  NAND2_X4 U3507 ( .A1(b[13]), .A2(a[13]), .ZN(net213443) );
  NAND2_X4 U3508 ( .A1(a[12]), .A2(b[12]), .ZN(net214022) );
  NAND2_X4 U3509 ( .A1(b[10]), .A2(a[10]), .ZN(net215210) );
  INV_X4 U3510 ( .A(net217237), .ZN(net220019) );
  NAND2_X1 U3511 ( .A1(net217235), .A2(net217082), .ZN(n3241) );
  NAND2_X2 U3512 ( .A1(n3239), .A2(n3240), .ZN(n3242) );
  NAND2_X2 U3513 ( .A1(n3241), .A2(n3242), .ZN(net217084) );
  INV_X4 U3514 ( .A(net217235), .ZN(n3239) );
  INV_X2 U3515 ( .A(net217082), .ZN(n3240) );
  INV_X4 U3516 ( .A(a[4]), .ZN(net219068) );
  NAND2_X2 U3517 ( .A1(net218626), .A2(a[4]), .ZN(n4418) );
  NAND2_X2 U3518 ( .A1(b[16]), .A2(a[4]), .ZN(net215301) );
  NAND2_X2 U3519 ( .A1(a[4]), .A2(b[27]), .ZN(n7688) );
  NAND2_X2 U3520 ( .A1(b[10]), .A2(a[4]), .ZN(n5204) );
  NAND2_X2 U3521 ( .A1(net218530), .A2(a[4]), .ZN(n4520) );
  AOI21_X2 U3522 ( .B1(n4594), .B2(net217442), .A(n4593), .ZN(n4595) );
  NOR2_X2 U3523 ( .A1(n4420), .A2(n4419), .ZN(n4422) );
  NAND3_X2 U3524 ( .A1(n4592), .A2(n4516), .A3(n4515), .ZN(n4603) );
  OAI21_X2 U3525 ( .B1(n4522), .B2(n4521), .A(n4592), .ZN(n4523) );
  NAND2_X2 U3526 ( .A1(a[3]), .A2(a[4]), .ZN(net219054) );
  INV_X8 U3527 ( .A(n6831), .ZN(n6962) );
  INV_X1 U3528 ( .A(net213223), .ZN(net213219) );
  INV_X8 U3529 ( .A(net212735), .ZN(net212732) );
  NAND2_X4 U3530 ( .A1(net213389), .A2(net213388), .ZN(n3243) );
  INV_X1 U3531 ( .A(net241088), .ZN(net241077) );
  NAND2_X2 U3532 ( .A1(n5628), .A2(n5630), .ZN(n5544) );
  NAND2_X4 U3533 ( .A1(net218240), .A2(net218257), .ZN(net218251) );
  NAND2_X4 U3534 ( .A1(n5833), .A2(n5834), .ZN(n5901) );
  NAND2_X4 U3535 ( .A1(n6148), .A2(n5894), .ZN(n5844) );
  NAND2_X4 U3536 ( .A1(n5840), .A2(n5841), .ZN(n6148) );
  NAND2_X4 U3537 ( .A1(net213019), .A2(net213384), .ZN(n3244) );
  NAND2_X2 U3538 ( .A1(n3243), .A2(net213384), .ZN(net212733) );
  INV_X4 U3539 ( .A(n5692), .ZN(n5691) );
  NAND2_X2 U3540 ( .A1(n6807), .A2(net213981), .ZN(n3247) );
  NAND2_X2 U3541 ( .A1(n3245), .A2(n3246), .ZN(n3248) );
  NAND2_X2 U3542 ( .A1(n3247), .A2(n3248), .ZN(n3874) );
  INV_X2 U3543 ( .A(n6807), .ZN(n3245) );
  INV_X4 U3544 ( .A(net213981), .ZN(n3246) );
  INV_X2 U3545 ( .A(net215105), .ZN(net215107) );
  INV_X1 U3546 ( .A(n7541), .ZN(n7545) );
  OAI21_X2 U3547 ( .B1(n7255), .B2(net212891), .A(n7254), .ZN(n7402) );
  INV_X4 U3548 ( .A(net212883), .ZN(net212881) );
  NAND3_X1 U3549 ( .A1(net212137), .A2(net212138), .A3(n3829), .ZN(n3828) );
  INV_X2 U3550 ( .A(net212137), .ZN(net212377) );
  NAND2_X1 U3551 ( .A1(n3344), .A2(n7765), .ZN(n7766) );
  CLKBUF_X3 U3552 ( .A(n7239), .Z(n3929) );
  INV_X2 U3553 ( .A(net212911), .ZN(net212909) );
  NAND2_X4 U3554 ( .A1(net213052), .A2(net220068), .ZN(net212924) );
  NAND2_X4 U3555 ( .A1(n6940), .A2(n3947), .ZN(net213707) );
  NAND2_X4 U3556 ( .A1(n3833), .A2(n3796), .ZN(net215342) );
  INV_X8 U3557 ( .A(net213598), .ZN(net213246) );
  INV_X4 U3558 ( .A(n6891), .ZN(n6894) );
  NAND2_X4 U3559 ( .A1(n3513), .A2(net213770), .ZN(net213551) );
  NAND2_X4 U3560 ( .A1(n7748), .A2(n7747), .ZN(n7511) );
  OAI211_X1 U3561 ( .C1(n3960), .C2(n3991), .A(net218608), .B(n3398), .ZN(
        n5738) );
  INV_X2 U3562 ( .A(n3960), .ZN(n5735) );
  XNOR2_X1 U3563 ( .A(n5864), .B(n5981), .ZN(n5867) );
  NAND2_X2 U3564 ( .A1(n5441), .A2(n5442), .ZN(net215476) );
  NAND2_X4 U3565 ( .A1(n3686), .A2(n3682), .ZN(net215447) );
  NAND2_X4 U3566 ( .A1(n6949), .A2(n6950), .ZN(n7113) );
  NAND2_X2 U3567 ( .A1(n5473), .A2(n5472), .ZN(n5637) );
  INV_X8 U3568 ( .A(n6896), .ZN(n6898) );
  INV_X2 U3569 ( .A(n4160), .ZN(n4158) );
  NAND2_X1 U3570 ( .A1(n5846), .A2(n5845), .ZN(n5890) );
  NAND2_X2 U3571 ( .A1(net214983), .A2(net215057), .ZN(n3703) );
  INV_X4 U3572 ( .A(n3670), .ZN(n3671) );
  INV_X2 U3573 ( .A(net213736), .ZN(net213578) );
  NAND2_X4 U3574 ( .A1(n3739), .A2(n3738), .ZN(n3736) );
  NAND2_X4 U3575 ( .A1(n3272), .A2(n4805), .ZN(n4806) );
  CLKBUF_X3 U3576 ( .A(n6939), .Z(n3947) );
  NAND2_X1 U3577 ( .A1(n5839), .A2(n5838), .ZN(n3251) );
  NAND2_X4 U3578 ( .A1(n3249), .A2(n3250), .ZN(n3252) );
  NAND2_X4 U3579 ( .A1(n3251), .A2(n3252), .ZN(n5841) );
  INV_X4 U3580 ( .A(n5839), .ZN(n3249) );
  INV_X4 U3581 ( .A(n5838), .ZN(n3250) );
  NAND2_X1 U3582 ( .A1(n3628), .A2(n3627), .ZN(n3255) );
  NAND2_X2 U3583 ( .A1(n3253), .A2(n3254), .ZN(n3256) );
  NAND2_X2 U3584 ( .A1(n3255), .A2(n3256), .ZN(net214795) );
  INV_X2 U3585 ( .A(n3628), .ZN(n3253) );
  INV_X2 U3586 ( .A(n3627), .ZN(n3254) );
  NAND2_X1 U3587 ( .A1(net215078), .A2(n3687), .ZN(n3258) );
  NAND2_X2 U3588 ( .A1(net215082), .A2(n3257), .ZN(n3259) );
  NAND2_X2 U3589 ( .A1(n3258), .A2(n3259), .ZN(net215075) );
  NAND2_X2 U3590 ( .A1(net214814), .A2(n3261), .ZN(n3262) );
  NAND2_X2 U3591 ( .A1(n3260), .A2(net214815), .ZN(n3263) );
  NAND2_X2 U3592 ( .A1(n3262), .A2(n3263), .ZN(net219429) );
  INV_X2 U3593 ( .A(net214814), .ZN(n3260) );
  INV_X4 U3594 ( .A(net214815), .ZN(n3261) );
  INV_X4 U3595 ( .A(n5841), .ZN(n5843) );
  NAND2_X4 U3596 ( .A1(net218269), .A2(net218217), .ZN(net218306) );
  INV_X8 U3597 ( .A(net214713), .ZN(net214711) );
  NAND2_X1 U3598 ( .A1(net212651), .A2(net212652), .ZN(net212650) );
  INV_X4 U3599 ( .A(net215812), .ZN(net215811) );
  NAND2_X4 U3600 ( .A1(net213809), .A2(net213524), .ZN(net213523) );
  NAND2_X4 U3601 ( .A1(net218576), .A2(a[9]), .ZN(net216885) );
  NAND2_X4 U3602 ( .A1(net218558), .A2(a[8]), .ZN(net217899) );
  NAND2_X2 U3603 ( .A1(net212389), .A2(net219445), .ZN(n3264) );
  INV_X2 U3604 ( .A(net212391), .ZN(n3265) );
  AND2_X2 U3605 ( .A1(n3264), .A2(n3265), .ZN(net212116) );
  NAND2_X2 U3606 ( .A1(net212113), .A2(net212112), .ZN(n3268) );
  NAND2_X4 U3607 ( .A1(n3266), .A2(n3267), .ZN(n3269) );
  NAND2_X4 U3608 ( .A1(n3268), .A2(n3269), .ZN(net212111) );
  INV_X4 U3609 ( .A(net212113), .ZN(n3266) );
  INV_X4 U3610 ( .A(net212112), .ZN(n3267) );
  NOR2_X4 U3611 ( .A1(net212392), .A2(net212393), .ZN(net212391) );
  NAND2_X1 U3612 ( .A1(net212399), .A2(net223009), .ZN(net212112) );
  NAND2_X4 U3613 ( .A1(a[3]), .A2(b[0]), .ZN(n3270) );
  NAND2_X4 U3614 ( .A1(n4051), .A2(n4050), .ZN(n4068) );
  INV_X2 U3615 ( .A(n4051), .ZN(n4049) );
  NAND2_X4 U3616 ( .A1(net218556), .A2(a[16]), .ZN(net215855) );
  NAND2_X4 U3617 ( .A1(n5639), .A2(n5638), .ZN(n5516) );
  INV_X2 U3618 ( .A(n4988), .ZN(n4895) );
  OR2_X2 U3619 ( .A1(n4987), .A2(n4895), .ZN(n3776) );
  OAI21_X2 U3620 ( .B1(n4895), .B2(n4894), .A(n4893), .ZN(n4898) );
  NAND2_X4 U3621 ( .A1(n6436), .A2(n6437), .ZN(n6674) );
  NAND2_X2 U3622 ( .A1(n3288), .A2(net218808), .ZN(net218809) );
  INV_X2 U3623 ( .A(n6089), .ZN(n6087) );
  INV_X1 U3624 ( .A(n4085), .ZN(n4088) );
  INV_X4 U3625 ( .A(net218136), .ZN(n3708) );
  NOR2_X4 U3626 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  OAI21_X4 U3627 ( .B1(n6677), .B2(n6676), .A(n6675), .ZN(n6606) );
  NAND2_X4 U3628 ( .A1(n5221), .A2(n5220), .ZN(n5255) );
  NAND2_X4 U3629 ( .A1(n5389), .A2(n5390), .ZN(n5638) );
  NAND2_X2 U3630 ( .A1(n4896), .A2(net216960), .ZN(n4897) );
  INV_X8 U3631 ( .A(n5649), .ZN(n5375) );
  INV_X4 U3632 ( .A(n5645), .ZN(n5646) );
  INV_X2 U3633 ( .A(n5507), .ZN(n3944) );
  INV_X2 U3634 ( .A(net213173), .ZN(net213169) );
  INV_X2 U3635 ( .A(net213132), .ZN(n3484) );
  NAND2_X4 U3636 ( .A1(net213130), .A2(net213132), .ZN(net213495) );
  NAND2_X4 U3637 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  NAND3_X4 U3638 ( .A1(net216190), .A2(net220521), .A3(net216191), .ZN(
        net215790) );
  INV_X8 U3639 ( .A(n5911), .ZN(n5912) );
  NAND2_X2 U3640 ( .A1(n4072), .A2(net218224), .ZN(net218219) );
  INV_X8 U3641 ( .A(n4087), .ZN(n4061) );
  NAND2_X4 U3642 ( .A1(n5097), .A2(n5232), .ZN(n5233) );
  INV_X1 U3643 ( .A(net212926), .ZN(net212922) );
  INV_X2 U3644 ( .A(n6172), .ZN(n6175) );
  NAND2_X4 U3645 ( .A1(n4046), .A2(net218091), .ZN(n4048) );
  NAND2_X2 U3646 ( .A1(n4119), .A2(net218091), .ZN(n3283) );
  INV_X2 U3647 ( .A(n4891), .ZN(n3271) );
  INV_X4 U3648 ( .A(n3271), .ZN(n3272) );
  NAND2_X1 U3649 ( .A1(n4904), .A2(n3274), .ZN(n3275) );
  NAND2_X2 U3650 ( .A1(n3273), .A2(n4903), .ZN(n3276) );
  NAND2_X2 U3651 ( .A1(n3275), .A2(n3276), .ZN(n3339) );
  INV_X1 U3652 ( .A(n4904), .ZN(n3273) );
  INV_X4 U3653 ( .A(n4903), .ZN(n3274) );
  NAND2_X2 U3654 ( .A1(n3277), .A2(n3278), .ZN(n3279) );
  NAND2_X4 U3655 ( .A1(n3279), .A2(n4979), .ZN(n4909) );
  INV_X4 U3656 ( .A(n3339), .ZN(n3277) );
  INV_X2 U3657 ( .A(n4971), .ZN(n3278) );
  NAND2_X4 U3658 ( .A1(b[4]), .A2(a[8]), .ZN(n4971) );
  NAND2_X4 U3659 ( .A1(n3742), .A2(net216767), .ZN(n3738) );
  NAND2_X4 U3660 ( .A1(n6399), .A2(n6400), .ZN(n6699) );
  NAND2_X4 U3661 ( .A1(net218576), .A2(a[6]), .ZN(n4050) );
  NAND2_X4 U3662 ( .A1(n6333), .A2(n6332), .ZN(n6533) );
  NAND2_X2 U3663 ( .A1(n5090), .A2(n3968), .ZN(n5360) );
  NAND2_X2 U3664 ( .A1(net217259), .A2(n4798), .ZN(n3280) );
  BUF_X8 U3665 ( .A(net215669), .Z(n3281) );
  INV_X2 U3666 ( .A(net218170), .ZN(net218096) );
  NAND2_X1 U3667 ( .A1(n5833), .A2(n5834), .ZN(n3282) );
  NAND2_X2 U3668 ( .A1(n3284), .A2(n4120), .ZN(n4047) );
  INV_X2 U3669 ( .A(n3283), .ZN(n3284) );
  INV_X2 U3670 ( .A(n5835), .ZN(n5833) );
  NAND2_X4 U3671 ( .A1(n4358), .A2(n4266), .ZN(net218091) );
  NAND2_X2 U3672 ( .A1(n3285), .A2(n3286), .ZN(n3287) );
  NAND2_X2 U3673 ( .A1(n3287), .A2(n5803), .ZN(n5804) );
  INV_X2 U3674 ( .A(n3307), .ZN(n3285) );
  INV_X4 U3675 ( .A(n3962), .ZN(n3286) );
  INV_X4 U3676 ( .A(n5804), .ZN(n5510) );
  NAND2_X4 U3677 ( .A1(net218576), .A2(a[10]), .ZN(net217271) );
  NAND2_X2 U3678 ( .A1(net218158), .A2(net218083), .ZN(net241366) );
  INV_X1 U3679 ( .A(n7538), .ZN(n7540) );
  NAND2_X2 U3680 ( .A1(net212390), .A2(net219412), .ZN(net212413) );
  NAND2_X1 U3681 ( .A1(n7580), .A2(n7579), .ZN(n7582) );
  INV_X8 U3682 ( .A(net214461), .ZN(net214808) );
  INV_X4 U3683 ( .A(n3838), .ZN(n3837) );
  NAND2_X4 U3684 ( .A1(n6806), .A2(n6805), .ZN(net213736) );
  OAI21_X4 U3685 ( .B1(net213870), .B2(net213560), .A(net213562), .ZN(n3481)
         );
  NAND2_X4 U3686 ( .A1(n4795), .A2(n4730), .ZN(n4129) );
  OAI21_X4 U3687 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5628) );
  NAND2_X4 U3688 ( .A1(n6419), .A2(n6420), .ZN(net213992) );
  NAND2_X2 U3689 ( .A1(net216839), .A2(net216578), .ZN(net217069) );
  XNOR2_X2 U3690 ( .A(net217082), .B(net216941), .ZN(net217081) );
  NAND2_X2 U3691 ( .A1(net216220), .A2(net216219), .ZN(net216217) );
  NAND2_X1 U3692 ( .A1(n6793), .A2(n6898), .ZN(n3291) );
  NAND2_X2 U3693 ( .A1(n3289), .A2(n3290), .ZN(n3292) );
  NAND2_X2 U3694 ( .A1(n3291), .A2(n3292), .ZN(n3873) );
  INV_X1 U3695 ( .A(n6898), .ZN(n3289) );
  NAND2_X4 U3696 ( .A1(net213737), .A2(n3293), .ZN(n3295) );
  INV_X4 U3697 ( .A(net213574), .ZN(n3293) );
  NAND2_X4 U3698 ( .A1(n3669), .A2(n3674), .ZN(net213587) );
  NAND2_X4 U3699 ( .A1(net218057), .A2(net217229), .ZN(net218133) );
  NAND2_X4 U3700 ( .A1(net223706), .A2(net219611), .ZN(n5818) );
  INV_X8 U3701 ( .A(net214818), .ZN(net214717) );
  NAND2_X4 U3702 ( .A1(n4753), .A2(n4752), .ZN(n4835) );
  NAND2_X4 U3703 ( .A1(n4823), .A2(n4829), .ZN(n4750) );
  INV_X4 U3704 ( .A(net215318), .ZN(net215320) );
  INV_X4 U3705 ( .A(net214719), .ZN(net214819) );
  NAND2_X4 U3706 ( .A1(net215107), .A2(net215106), .ZN(n3624) );
  INV_X2 U3707 ( .A(net218267), .ZN(net218260) );
  NAND2_X4 U3708 ( .A1(b[4]), .A2(a[4]), .ZN(net217244) );
  NOR2_X4 U3709 ( .A1(n3297), .A2(n3298), .ZN(n3296) );
  INV_X32 U3710 ( .A(a[3]), .ZN(n3297) );
  INV_X4 U3711 ( .A(n4901), .ZN(n4899) );
  NAND2_X4 U3712 ( .A1(n5895), .A2(n5891), .ZN(n5709) );
  NAND2_X4 U3713 ( .A1(b[0]), .A2(a[2]), .ZN(n3881) );
  NAND2_X4 U3714 ( .A1(b[0]), .A2(a[5]), .ZN(n3910) );
  NAND2_X4 U3715 ( .A1(b[0]), .A2(a[2]), .ZN(n3880) );
  NAND2_X4 U3716 ( .A1(b[0]), .A2(a[5]), .ZN(n3909) );
  NAND2_X4 U3717 ( .A1(b[0]), .A2(a[5]), .ZN(n4484) );
  NAND2_X4 U3718 ( .A1(b[1]), .A2(b[0]), .ZN(net220395) );
  INV_X4 U3719 ( .A(n6707), .ZN(n6498) );
  CLKBUF_X2 U3720 ( .A(net216841), .Z(n3299) );
  INV_X8 U3721 ( .A(net216285), .ZN(net216281) );
  NAND2_X4 U3722 ( .A1(n6564), .A2(n6565), .ZN(n6722) );
  NAND2_X4 U3723 ( .A1(n6032), .A2(n6031), .ZN(n6163) );
  OAI21_X4 U3724 ( .B1(n5370), .B2(n5491), .A(n5496), .ZN(n5372) );
  XNOR2_X2 U3725 ( .A(net216768), .B(net216769), .ZN(net216767) );
  INV_X4 U3726 ( .A(net215061), .ZN(n3702) );
  NAND2_X2 U3727 ( .A1(net215064), .A2(n6085), .ZN(n3582) );
  INV_X4 U3728 ( .A(n4791), .ZN(n4882) );
  INV_X8 U3729 ( .A(net218114), .ZN(net217237) );
  NAND2_X4 U3730 ( .A1(net218076), .A2(n4123), .ZN(net217259) );
  NOR2_X4 U3731 ( .A1(n3570), .A2(n3646), .ZN(n3649) );
  XNOR2_X2 U3732 ( .A(n3173), .B(n5354), .ZN(n5252) );
  INV_X8 U3733 ( .A(net217290), .ZN(net219864) );
  NOR2_X4 U3734 ( .A1(net218161), .A2(n3301), .ZN(n3300) );
  INV_X4 U3735 ( .A(n3300), .ZN(net217028) );
  INV_X4 U3736 ( .A(net218161), .ZN(net217970) );
  NAND2_X4 U3737 ( .A1(n6194), .A2(n6195), .ZN(n6322) );
  INV_X2 U3738 ( .A(net218245), .ZN(net218262) );
  NAND2_X4 U3739 ( .A1(n4092), .A2(net218115), .ZN(n4108) );
  AOI21_X4 U3740 ( .B1(n4800), .B2(net216811), .A(n4989), .ZN(n4801) );
  NAND2_X4 U3741 ( .A1(n6558), .A2(n6559), .ZN(n6728) );
  NAND2_X4 U3742 ( .A1(n7368), .A2(n3898), .ZN(n7551) );
  NAND2_X4 U3743 ( .A1(n7314), .A2(n7315), .ZN(n7403) );
  NAND2_X4 U3744 ( .A1(n7337), .A2(n3200), .ZN(n7514) );
  OAI21_X4 U3745 ( .B1(net212871), .B2(n7267), .A(n7266), .ZN(n7424) );
  NAND2_X4 U3746 ( .A1(net216644), .A2(net216285), .ZN(n5219) );
  NAND2_X4 U3747 ( .A1(net218219), .A2(net218220), .ZN(net218173) );
  CLKBUF_X3 U3748 ( .A(n5803), .Z(n3572) );
  NAND2_X1 U3749 ( .A1(n6682), .A2(n6878), .ZN(n6599) );
  NAND2_X4 U3750 ( .A1(n4040), .A2(n4039), .ZN(net218266) );
  XNOR2_X2 U3751 ( .A(net220397), .B(n4038), .ZN(n4039) );
  NAND2_X4 U3752 ( .A1(net213491), .A2(net213492), .ZN(net213168) );
  XNOR2_X1 U3753 ( .A(n4033), .B(n4035), .ZN(n4030) );
  INV_X4 U3754 ( .A(n7184), .ZN(n7182) );
  INV_X4 U3755 ( .A(n6305), .ZN(n6306) );
  INV_X4 U3756 ( .A(net213758), .ZN(n3817) );
  NAND2_X4 U3757 ( .A1(net216092), .A2(net215797), .ZN(n3651) );
  INV_X8 U3758 ( .A(net214619), .ZN(net214427) );
  NAND2_X4 U3759 ( .A1(n5488), .A2(net216063), .ZN(n5783) );
  INV_X4 U3760 ( .A(n3302), .ZN(net220017) );
  NAND2_X4 U3761 ( .A1(net213221), .A2(net213223), .ZN(net213419) );
  NAND2_X2 U3762 ( .A1(n6383), .A2(n6382), .ZN(n3591) );
  INV_X4 U3763 ( .A(net213597), .ZN(n3302) );
  INV_X4 U3764 ( .A(net213597), .ZN(net213247) );
  NAND4_X1 U3765 ( .A1(n5045), .A2(n5044), .A3(net216710), .A4(net216711), 
        .ZN(n6850) );
  AND4_X2 U3766 ( .A1(net217029), .A2(n5044), .A3(net217816), .A4(n4447), .ZN(
        n3333) );
  INV_X4 U3767 ( .A(n6712), .ZN(n6509) );
  NAND2_X4 U3768 ( .A1(n5931), .A2(n6044), .ZN(n6045) );
  INV_X2 U3769 ( .A(n5930), .ZN(n5928) );
  NAND2_X1 U3770 ( .A1(n3445), .A2(net217271), .ZN(n3444) );
  NAND2_X4 U3771 ( .A1(n3897), .A2(n5547), .ZN(n5904) );
  NAND2_X4 U3772 ( .A1(n6090), .A2(n6089), .ZN(n6426) );
  NAND2_X4 U3773 ( .A1(net219236), .A2(net219237), .ZN(n3696) );
  INV_X8 U3774 ( .A(n5479), .ZN(n5805) );
  NAND2_X4 U3775 ( .A1(net216653), .A2(net217228), .ZN(n4728) );
  NAND2_X4 U3776 ( .A1(n5473), .A2(n5471), .ZN(n5283) );
  NAND2_X4 U3777 ( .A1(n4728), .A2(n4727), .ZN(n4794) );
  INV_X4 U3778 ( .A(n4986), .ZN(n4992) );
  INV_X8 U3779 ( .A(net216282), .ZN(net216644) );
  NAND2_X2 U3780 ( .A1(n6221), .A2(net214603), .ZN(n3800) );
  NAND2_X4 U3781 ( .A1(net213570), .A2(net213572), .ZN(n3536) );
  NAND2_X2 U3782 ( .A1(n6313), .A2(n6310), .ZN(n6210) );
  INV_X4 U3783 ( .A(net214543), .ZN(net214541) );
  INV_X2 U3784 ( .A(net214714), .ZN(net214710) );
  INV_X2 U3785 ( .A(n4067), .ZN(n4266) );
  INV_X4 U3786 ( .A(n5091), .ZN(n5242) );
  INV_X8 U3787 ( .A(n5243), .ZN(n5361) );
  NAND2_X4 U3788 ( .A1(n5241), .A2(n5242), .ZN(n5243) );
  NAND2_X4 U3789 ( .A1(net214713), .A2(n3588), .ZN(net214840) );
  NAND2_X4 U3790 ( .A1(n5771), .A2(n3605), .ZN(n5681) );
  NOR2_X2 U3791 ( .A1(net219162), .A2(n3635), .ZN(n3629) );
  NAND2_X4 U3792 ( .A1(n3679), .A2(net215569), .ZN(net215215) );
  OAI211_X4 U3793 ( .C1(net216281), .C2(net216282), .A(net216283), .B(
        net216284), .ZN(net216279) );
  XNOR2_X2 U3794 ( .A(net213576), .B(net213997), .ZN(n3503) );
  NAND2_X2 U3795 ( .A1(n6901), .A2(n6900), .ZN(n6904) );
  OAI21_X2 U3796 ( .B1(n6523), .B2(n6522), .A(n6521), .ZN(n6525) );
  NOR2_X4 U3797 ( .A1(net217140), .A2(net217141), .ZN(net217127) );
  NAND2_X2 U3798 ( .A1(n5918), .A2(n6035), .ZN(n6036) );
  NAND2_X4 U3799 ( .A1(n7505), .A2(n7502), .ZN(n7335) );
  NAND2_X4 U3800 ( .A1(n7257), .A2(n7256), .ZN(n7156) );
  NAND2_X4 U3801 ( .A1(net215186), .A2(net215185), .ZN(net215417) );
  NAND2_X4 U3802 ( .A1(n6348), .A2(n6537), .ZN(n6538) );
  INV_X16 U3803 ( .A(n7855), .ZN(n3999) );
  NAND2_X2 U3804 ( .A1(n7131), .A2(n7266), .ZN(n7267) );
  NOR2_X2 U3805 ( .A1(net217545), .A2(n4509), .ZN(n4511) );
  NOR2_X1 U3806 ( .A1(net218556), .A2(net218484), .ZN(n4510) );
  NOR2_X2 U3807 ( .A1(net217529), .A2(n4520), .ZN(n4522) );
  OAI21_X2 U3808 ( .B1(n4600), .B2(n4599), .A(net217431), .ZN(n4602) );
  OAI21_X2 U3809 ( .B1(n4576), .B2(n4543), .A(n4542), .ZN(n4545) );
  NOR2_X2 U3810 ( .A1(b[16]), .A2(net216124), .ZN(n4544) );
  NOR2_X1 U3811 ( .A1(n4550), .A2(n5998), .ZN(n4552) );
  NOR2_X2 U3812 ( .A1(b[18]), .A2(net215709), .ZN(n4549) );
  NOR2_X2 U3813 ( .A1(b[19]), .A2(net215499), .ZN(n4548) );
  OAI21_X2 U3814 ( .B1(n4565), .B2(n7001), .A(n4564), .ZN(n4567) );
  NOR3_X2 U3815 ( .A1(n4585), .A2(n4584), .A3(n4583), .ZN(n4586) );
  INV_X4 U3816 ( .A(n7871), .ZN(n3994) );
  NOR2_X2 U3817 ( .A1(op[0]), .A2(n3457), .ZN(net217960) );
  OAI21_X2 U3818 ( .B1(n4269), .B2(n4268), .A(n7039), .ZN(n4270) );
  NOR2_X1 U3819 ( .A1(n5058), .A2(n3996), .ZN(n4394) );
  NOR2_X1 U3820 ( .A1(n5181), .A2(n3996), .ZN(n4428) );
  NOR2_X1 U3821 ( .A1(net216306), .A2(n3996), .ZN(n4461) );
  INV_X4 U3822 ( .A(net218542), .ZN(net218540) );
  OAI21_X2 U3823 ( .B1(n3340), .B2(n7460), .A(n7711), .ZN(n7463) );
  NAND2_X2 U3824 ( .A1(n3324), .A2(n7290), .ZN(n7420) );
  NAND2_X2 U3825 ( .A1(net213542), .A2(net213543), .ZN(net213779) );
  INV_X4 U3826 ( .A(net214569), .ZN(net215081) );
  INV_X4 U3827 ( .A(net215091), .ZN(net215087) );
  NAND2_X2 U3828 ( .A1(n5216), .A2(net216202), .ZN(n5124) );
  AOI211_X2 U3829 ( .C1(n4608), .C2(n4607), .A(n4606), .B(n4605), .ZN(n4611)
         );
  OAI21_X1 U3830 ( .B1(n4525), .B2(n4524), .A(n4607), .ZN(n4527) );
  AOI21_X2 U3831 ( .B1(n5554), .B2(n5627), .A(n5553), .ZN(n5555) );
  NOR2_X2 U3832 ( .A1(a[19]), .A2(net217395), .ZN(n4627) );
  INV_X4 U3833 ( .A(n3528), .ZN(n3527) );
  OAI21_X2 U3834 ( .B1(n4547), .B2(n5605), .A(n4546), .ZN(n4557) );
  AOI21_X2 U3835 ( .B1(n4554), .B2(n4553), .A(n4635), .ZN(n4555) );
  OAI21_X2 U3836 ( .B1(n4552), .B2(n4551), .A(n6108), .ZN(n4553) );
  NOR2_X2 U3837 ( .A1(b[20]), .A2(net215252), .ZN(n4551) );
  NOR2_X2 U3838 ( .A1(b[22]), .A2(net214758), .ZN(n4556) );
  OAI21_X2 U3839 ( .B1(n4569), .B2(n4653), .A(n4568), .ZN(n4571) );
  NOR2_X2 U3840 ( .A1(b[27]), .A2(n7054), .ZN(n4566) );
  NOR2_X2 U3841 ( .A1(b[29]), .A2(n7387), .ZN(n4570) );
  NOR3_X1 U3842 ( .A1(n4658), .A2(n4610), .A3(n4642), .ZN(n4589) );
  NOR3_X1 U3843 ( .A1(n4576), .A2(n4603), .A3(n4591), .ZN(n4588) );
  NAND3_X2 U3844 ( .A1(b[8]), .A2(a[0]), .A3(n4477), .ZN(n4824) );
  NAND3_X2 U3845 ( .A1(b[12]), .A2(a[0]), .A3(n5033), .ZN(n5150) );
  NAND3_X2 U3846 ( .A1(b[13]), .A2(a[0]), .A3(n5157), .ZN(n5197) );
  NAND3_X2 U3847 ( .A1(b[14]), .A2(a[0]), .A3(n5306), .ZN(n5568) );
  NAND3_X2 U3848 ( .A1(b[25]), .A2(a[0]), .A3(n6972), .ZN(n7105) );
  NOR2_X1 U3849 ( .A1(n7223), .A2(n3995), .ZN(n7224) );
  NOR2_X1 U3850 ( .A1(net212005), .A2(n3993), .ZN(n7874) );
  NOR2_X1 U3851 ( .A1(net212008), .A2(n7869), .ZN(n7875) );
  NOR2_X2 U3852 ( .A1(n7872), .A2(n3995), .ZN(n7873) );
  OAI21_X1 U3853 ( .B1(n4682), .B2(n3995), .A(n4681), .ZN(n4683) );
  NOR2_X1 U3854 ( .A1(n4943), .A2(n7869), .ZN(n4684) );
  NAND3_X2 U3855 ( .A1(n4221), .A2(n4220), .A3(n4219), .ZN(n4241) );
  NOR2_X1 U3856 ( .A1(net218554), .A2(n3991), .ZN(net217877) );
  INV_X4 U3857 ( .A(a[1]), .ZN(net218486) );
  NOR2_X1 U3858 ( .A1(n3360), .A2(n5332), .ZN(n4395) );
  NAND2_X2 U3859 ( .A1(n4085), .A2(n4086), .ZN(n4081) );
  NOR2_X1 U3860 ( .A1(n4777), .A2(n5332), .ZN(n4429) );
  NOR2_X1 U3861 ( .A1(n4460), .A2(n5332), .ZN(n4462) );
  INV_X16 U3862 ( .A(net218658), .ZN(net218659) );
  AOI21_X2 U3863 ( .B1(n7803), .B2(n5595), .A(n5043), .ZN(n5047) );
  NOR2_X1 U3864 ( .A1(n5042), .A2(n7869), .ZN(n5043) );
  INV_X16 U3865 ( .A(n3377), .ZN(n3996) );
  OAI21_X1 U3866 ( .B1(net218544), .B2(n7038), .A(n4320), .ZN(n4319) );
  NAND3_X2 U3867 ( .A1(n4344), .A2(n4343), .A3(n4342), .ZN(n6005) );
  OAI21_X1 U3868 ( .B1(n3995), .B2(n7863), .A(n4452), .ZN(n6467) );
  NOR2_X1 U3869 ( .A1(n7081), .A2(n7079), .ZN(n6635) );
  NOR2_X1 U3870 ( .A1(n6645), .A2(n3332), .ZN(n6647) );
  NOR2_X1 U3871 ( .A1(n6001), .A2(n3373), .ZN(n6003) );
  OAI21_X1 U3872 ( .B1(n4193), .B2(n3993), .A(n4192), .ZN(n4194) );
  AOI21_X2 U3873 ( .B1(n7805), .B2(n7831), .A(n4773), .ZN(n6977) );
  NOR2_X1 U3874 ( .A1(net212677), .A2(n7378), .ZN(net212673) );
  NOR2_X1 U3875 ( .A1(b[29]), .A2(net218660), .ZN(n7378) );
  NOR2_X1 U3876 ( .A1(n7889), .A2(net218606), .ZN(n7826) );
  NOR2_X1 U3877 ( .A1(net218496), .A2(n3460), .ZN(net212105) );
  INV_X8 U3878 ( .A(n3991), .ZN(n5193) );
  NOR2_X1 U3879 ( .A1(net218660), .A2(n4677), .ZN(n4275) );
  NOR2_X1 U3880 ( .A1(net218484), .A2(net218606), .ZN(n4262) );
  NAND3_X1 U3881 ( .A1(n4387), .A2(n4416), .A3(n4386), .ZN(n6113) );
  NOR2_X1 U3882 ( .A1(n6633), .A2(n6983), .ZN(n5447) );
  OAI21_X1 U3883 ( .B1(n5592), .B2(n5591), .A(n7036), .ZN(n5593) );
  NOR2_X2 U3884 ( .A1(net212677), .A2(n5590), .ZN(n5591) );
  NOR2_X2 U3885 ( .A1(b[17]), .A2(net218660), .ZN(n5590) );
  OAI21_X1 U3886 ( .B1(n5607), .B2(n6637), .A(n5606), .ZN(n5608) );
  NOR2_X1 U3887 ( .A1(net218378), .A2(net218608), .ZN(n5609) );
  NOR2_X2 U3888 ( .A1(b[18]), .A2(net218660), .ZN(n5733) );
  OAI21_X1 U3889 ( .B1(n5867), .B2(n5866), .A(n7036), .ZN(n5869) );
  NOR2_X2 U3890 ( .A1(net212677), .A2(n5865), .ZN(n5866) );
  NOR2_X2 U3891 ( .A1(b[19]), .A2(net218660), .ZN(n5865) );
  NOR2_X1 U3892 ( .A1(n6453), .A2(n6454), .ZN(n5868) );
  NOR2_X2 U3893 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NOR2_X2 U3894 ( .A1(net212677), .A2(n5986), .ZN(n5987) );
  NOR2_X2 U3895 ( .A1(b[20]), .A2(net218660), .ZN(n5986) );
  OAI21_X1 U3896 ( .B1(n7078), .B2(n3381), .A(n7036), .ZN(n5990) );
  OAI21_X1 U3897 ( .B1(n3369), .B2(n6637), .A(n6006), .ZN(n6007) );
  AOI21_X1 U3898 ( .B1(n6468), .B2(n6005), .A(n6004), .ZN(n6006) );
  NOR2_X1 U3899 ( .A1(n3364), .A2(n6135), .ZN(n6004) );
  NOR2_X1 U3900 ( .A1(n7081), .A2(n6983), .ZN(n5993) );
  NOR2_X1 U3901 ( .A1(n7074), .A2(n7053), .ZN(n5994) );
  NOR2_X1 U3902 ( .A1(n7080), .A2(n6984), .ZN(n5992) );
  NOR2_X1 U3903 ( .A1(n6124), .A2(n6983), .ZN(n6125) );
  NOR2_X1 U3904 ( .A1(n6122), .A2(n6984), .ZN(n6126) );
  AOI21_X1 U3905 ( .B1(n6099), .B2(net212094), .A(n6121), .ZN(n6104) );
  NOR2_X1 U3906 ( .A1(net214476), .A2(n6983), .ZN(n6477) );
  NOR2_X1 U3907 ( .A1(net214478), .A2(n6984), .ZN(n6478) );
  AOI21_X2 U3908 ( .B1(n6450), .B2(net212094), .A(n6449), .ZN(n6457) );
  OAI21_X1 U3909 ( .B1(n6844), .B2(n6843), .A(n7036), .ZN(n6847) );
  NOR2_X1 U3910 ( .A1(net212677), .A2(n6842), .ZN(n6843) );
  NOR2_X1 U3911 ( .A1(b[25]), .A2(net218660), .ZN(n6842) );
  NOR2_X1 U3912 ( .A1(n6845), .A2(n7035), .ZN(n6846) );
  OAI21_X1 U3913 ( .B1(n6861), .B2(n7058), .A(n6860), .ZN(n6862) );
  NOR2_X1 U3914 ( .A1(net213919), .A2(net218608), .ZN(n6863) );
  INV_X8 U3915 ( .A(n7053), .ZN(n6851) );
  OAI21_X1 U3916 ( .B1(n6976), .B2(n6975), .A(n7036), .ZN(n6979) );
  NOR2_X1 U3917 ( .A1(net212677), .A2(n6974), .ZN(n6975) );
  NOR2_X1 U3918 ( .A1(b[26]), .A2(net218660), .ZN(n6974) );
  NOR2_X1 U3919 ( .A1(n6977), .A2(n7035), .ZN(n6978) );
  OAI21_X1 U3920 ( .B1(n7003), .B2(n7058), .A(n7002), .ZN(n7004) );
  NOR2_X1 U3921 ( .A1(n6999), .A2(net218608), .ZN(n7005) );
  NOR2_X1 U3922 ( .A1(n6277), .A2(n6983), .ZN(n6987) );
  NOR2_X1 U3923 ( .A1(n6981), .A2(n7053), .ZN(n6988) );
  NOR2_X1 U3924 ( .A1(n6985), .A2(n6984), .ZN(n6986) );
  OAI21_X1 U3925 ( .B1(n7038), .B2(n3380), .A(net212061), .ZN(n7043) );
  NOR2_X1 U3926 ( .A1(n7041), .A2(n7828), .ZN(n7042) );
  OAI21_X1 U3927 ( .B1(n7059), .B2(n7058), .A(n7057), .ZN(n7060) );
  NOR2_X1 U3928 ( .A1(n7054), .A2(net218608), .ZN(n7061) );
  AOI21_X1 U3929 ( .B1(n7071), .B2(n7070), .A(n7818), .ZN(n7072) );
  AOI21_X2 U3930 ( .B1(n7208), .B2(net212094), .A(n7207), .ZN(n7209) );
  AOI21_X1 U3931 ( .B1(n7820), .B2(n7819), .A(n7818), .ZN(n7822) );
  OAI21_X1 U3932 ( .B1(n7889), .B2(net218600), .A(net218610), .ZN(n7890) );
  NAND3_X2 U3933 ( .A1(op[2]), .A2(n3455), .A3(net217346), .ZN(n3158) );
  OAI21_X2 U3934 ( .B1(net215177), .B2(net215178), .A(net214930), .ZN(
        net215175) );
  AOI21_X2 U3935 ( .B1(n5946), .B2(n5945), .A(n5944), .ZN(n5951) );
  OAI21_X2 U3936 ( .B1(net214662), .B2(net214663), .A(net214395), .ZN(
        net214660) );
  AOI21_X2 U3937 ( .B1(net214958), .B2(net223455), .A(net214959), .ZN(
        net214955) );
  OAI21_X2 U3938 ( .B1(n7015), .B2(net213508), .A(n7114), .ZN(n7017) );
  NAND2_X2 U3939 ( .A1(net213527), .A2(net213529), .ZN(n3548) );
  OAI21_X2 U3940 ( .B1(n5244), .B2(n5360), .A(n5359), .ZN(n5245) );
  INV_X4 U3941 ( .A(net215663), .ZN(n3612) );
  INV_X4 U3942 ( .A(n7265), .ZN(n7136) );
  OAI21_X1 U3943 ( .B1(n7434), .B2(n7817), .A(n7433), .ZN(n7637) );
  AOI21_X2 U3944 ( .B1(n7631), .B2(n7630), .A(n7629), .ZN(n7708) );
  INV_X4 U3945 ( .A(net216393), .ZN(net216221) );
  INV_X4 U3946 ( .A(n6017), .ZN(n6018) );
  OAI21_X2 U3947 ( .B1(n7626), .B2(n7625), .A(n7624), .ZN(n7714) );
  NAND2_X2 U3948 ( .A1(net214972), .A2(net214971), .ZN(net215096) );
  AOI21_X2 U3949 ( .B1(n7618), .B2(n7617), .A(n7616), .ZN(n7720) );
  OAI21_X2 U3950 ( .B1(n7611), .B2(n7610), .A(n7609), .ZN(n7726) );
  INV_X4 U3951 ( .A(n6246), .ZN(n3981) );
  NAND2_X2 U3952 ( .A1(n5350), .A2(n5525), .ZN(n5399) );
  AOI21_X1 U3953 ( .B1(net217433), .B2(net218496), .A(n4598), .ZN(n4599) );
  INV_X4 U3954 ( .A(n3602), .ZN(net219540) );
  OAI21_X1 U3955 ( .B1(n4595), .B2(net217438), .A(net217439), .ZN(n4596) );
  OAI21_X2 U3956 ( .B1(n4511), .B2(n4510), .A(n4582), .ZN(n4512) );
  AOI21_X2 U3957 ( .B1(net217524), .B2(n4523), .A(net217526), .ZN(n4525) );
  OAI21_X2 U3958 ( .B1(n6677), .B2(n6676), .A(n6675), .ZN(n6679) );
  NOR3_X2 U3959 ( .A1(b[9]), .A2(net217517), .A3(net218428), .ZN(n4529) );
  NOR2_X2 U3960 ( .A1(n4137), .A2(n4135), .ZN(n4115) );
  NAND2_X2 U3961 ( .A1(n3538), .A2(n3537), .ZN(net212454) );
  AOI21_X2 U3962 ( .B1(n5291), .B2(n5290), .A(n3870), .ZN(n5293) );
  AOI21_X1 U3963 ( .B1(n6108), .B2(n4632), .A(n4631), .ZN(n4636) );
  NOR2_X1 U3964 ( .A1(a[21]), .A2(net215232), .ZN(n4631) );
  OAI21_X1 U3965 ( .B1(n4630), .B2(n5998), .A(n4629), .ZN(n4632) );
  OAI21_X1 U3966 ( .B1(n4625), .B2(n5453), .A(n4624), .ZN(n4639) );
  AOI21_X1 U3967 ( .B1(n4622), .B2(n5190), .A(n4621), .ZN(n4625) );
  NOR2_X2 U3968 ( .A1(a[15]), .A2(net217403), .ZN(n4621) );
  NAND2_X2 U3969 ( .A1(n5208), .A2(n5212), .ZN(n5138) );
  INV_X4 U3970 ( .A(n5846), .ZN(n5614) );
  NOR2_X2 U3971 ( .A1(n7576), .A2(n7575), .ZN(n7577) );
  AOI211_X2 U3972 ( .C1(n4640), .C2(n4639), .A(n4638), .B(n4637), .ZN(n4643)
         );
  NOR2_X2 U3973 ( .A1(a[22]), .A2(net214984), .ZN(n4637) );
  NOR2_X1 U3974 ( .A1(n5605), .A2(n4591), .ZN(n4640) );
  OAI21_X2 U3975 ( .B1(n4636), .B2(n4635), .A(n4634), .ZN(n4638) );
  INV_X4 U3976 ( .A(n4026), .ZN(n4021) );
  AOI211_X2 U3977 ( .C1(n4633), .C2(n4557), .A(n4556), .B(n4555), .ZN(n4559)
         );
  NOR2_X2 U3978 ( .A1(b[25]), .A2(net213919), .ZN(n4561) );
  NOR2_X1 U3979 ( .A1(n6859), .A2(n7001), .ZN(n4578) );
  AOI21_X2 U3980 ( .B1(n3329), .B2(net217244), .A(net217529), .ZN(n4516) );
  NAND2_X2 U3981 ( .A1(n6297), .A2(n6291), .ZN(n6264) );
  OAI22_X2 U3982 ( .A1(n3766), .A2(n7234), .B1(n7026), .B2(n3926), .ZN(n7027)
         );
  NOR2_X2 U3983 ( .A1(n3460), .A2(net217356), .ZN(net217360) );
  AOI21_X2 U3984 ( .B1(n7230), .B2(n4571), .A(n4570), .ZN(n4573) );
  OAI21_X1 U3985 ( .B1(net217732), .B2(net218640), .A(net218610), .ZN(n4352)
         );
  NOR2_X1 U3986 ( .A1(n4334), .A2(n7069), .ZN(n7070) );
  NOR3_X2 U3987 ( .A1(n7084), .A2(n7083), .A3(n7082), .ZN(n7085) );
  NOR2_X1 U3988 ( .A1(n7080), .A2(n7079), .ZN(n7083) );
  NOR2_X1 U3989 ( .A1(n7081), .A2(n3993), .ZN(n7082) );
  NOR2_X1 U3990 ( .A1(net218544), .A2(n7078), .ZN(n7084) );
  NOR2_X2 U3991 ( .A1(n7077), .A2(n7076), .ZN(n7086) );
  NOR2_X1 U3992 ( .A1(n3364), .A2(n3995), .ZN(n7077) );
  NOR2_X1 U3993 ( .A1(n7387), .A2(net218600), .ZN(n7376) );
  NOR2_X1 U3994 ( .A1(net218558), .A2(n7217), .ZN(n7218) );
  NOR3_X2 U3995 ( .A1(n7226), .A2(n7225), .A3(n7224), .ZN(n7227) );
  NOR2_X1 U3996 ( .A1(net212970), .A2(n3993), .ZN(n7225) );
  NOR2_X1 U3997 ( .A1(n7221), .A2(n7869), .ZN(n7226) );
  AOI21_X2 U3998 ( .B1(n7851), .B2(n7850), .A(n7849), .ZN(n7853) );
  NOR2_X1 U3999 ( .A1(n7848), .A2(n7889), .ZN(n7849) );
  OAI21_X2 U4000 ( .B1(n7868), .B2(n7867), .A(n7866), .ZN(n7880) );
  NOR2_X1 U4001 ( .A1(net211993), .A2(net218640), .ZN(n7881) );
  NOR2_X1 U4002 ( .A1(net212023), .A2(net218600), .ZN(n7857) );
  NOR2_X1 U4003 ( .A1(n4668), .A2(net217346), .ZN(n4669) );
  OAI21_X2 U4004 ( .B1(n4679), .B2(n4678), .A(n7866), .ZN(n4694) );
  AOI21_X2 U4005 ( .B1(n4702), .B2(net218610), .A(n4701), .ZN(n4703) );
  NOR2_X1 U4006 ( .A1(net218600), .A2(n4700), .ZN(n4503) );
  NOR2_X1 U4007 ( .A1(n4207), .A2(n4942), .ZN(n4208) );
  NOR2_X2 U4008 ( .A1(n4206), .A2(n4205), .ZN(n4207) );
  NOR2_X2 U4009 ( .A1(n4779), .A2(n3996), .ZN(n4240) );
  AOI21_X2 U4010 ( .B1(n4237), .B2(n4236), .A(n6653), .ZN(n4238) );
  NOR2_X2 U4011 ( .A1(n4244), .A2(net218606), .ZN(n4239) );
  NOR2_X1 U4012 ( .A1(n4248), .A2(net218598), .ZN(n4250) );
  NOR2_X1 U4013 ( .A1(net218544), .A2(n7888), .ZN(n4309) );
  OAI21_X2 U4014 ( .B1(n5880), .B2(n4860), .A(n4321), .ZN(n4322) );
  NOR2_X1 U4015 ( .A1(n6453), .A2(n6135), .ZN(n4323) );
  NOR2_X2 U4016 ( .A1(b[4]), .A2(net218659), .ZN(n4327) );
  NOR2_X1 U4017 ( .A1(n4362), .A2(n4942), .ZN(n4371) );
  NOR2_X1 U4018 ( .A1(n4345), .A2(n4860), .ZN(n4346) );
  OAI21_X1 U4019 ( .B1(net217677), .B2(n4942), .A(n4398), .ZN(n4399) );
  AOI21_X2 U4020 ( .B1(n4775), .B2(net216704), .A(n4393), .ZN(n4397) );
  NOR2_X1 U4021 ( .A1(n4392), .A2(net218606), .ZN(n4393) );
  NOR2_X1 U4022 ( .A1(n6102), .A2(n6135), .ZN(n4388) );
  NOR2_X1 U4023 ( .A1(net217083), .A2(net218598), .ZN(n4377) );
  NOR2_X1 U4024 ( .A1(net218640), .A2(net217445), .ZN(n4378) );
  NOR2_X2 U4025 ( .A1(net212677), .A2(n4379), .ZN(n4381) );
  NOR2_X2 U4026 ( .A1(b[5]), .A2(net218659), .ZN(n4379) );
  OAI21_X1 U4027 ( .B1(n4434), .B2(n4942), .A(n4433), .ZN(n4435) );
  AOI21_X1 U4028 ( .B1(n4775), .B2(n5167), .A(n4426), .ZN(n4431) );
  NOR2_X1 U4029 ( .A1(n4425), .A2(net218606), .ZN(n4426) );
  NOR2_X1 U4030 ( .A1(n6273), .A2(n6135), .ZN(n4423) );
  NAND3_X1 U4031 ( .A1(n4417), .A2(n4416), .A3(n4415), .ZN(n6131) );
  NOR2_X1 U4032 ( .A1(net218640), .A2(n4592), .ZN(n4408) );
  NOR2_X1 U4033 ( .A1(net216979), .A2(net218598), .ZN(n4407) );
  NOR2_X2 U4034 ( .A1(net212677), .A2(n4409), .ZN(n4413) );
  OAI21_X1 U4035 ( .B1(n3333), .B2(n4942), .A(n4465), .ZN(n4466) );
  AOI21_X1 U4036 ( .B1(n4775), .B2(n5320), .A(n4459), .ZN(n4464) );
  NOR2_X1 U4037 ( .A1(net217608), .A2(net218606), .ZN(n4459) );
  NOR2_X1 U4038 ( .A1(n4453), .A2(n4768), .ZN(n4454) );
  NOR2_X1 U4039 ( .A1(n4451), .A2(n4860), .ZN(n4455) );
  NOR2_X1 U4040 ( .A1(net216394), .A2(net218598), .ZN(net217630) );
  NOR2_X1 U4041 ( .A1(net218640), .A2(net217439), .ZN(n4442) );
  NOR2_X2 U4042 ( .A1(net212677), .A2(n4443), .ZN(n4445) );
  NOR2_X2 U4043 ( .A1(b[7]), .A2(net218659), .ZN(n4443) );
  OAI21_X1 U4044 ( .B1(n7081), .B2(n6135), .A(n4488), .ZN(n4490) );
  NOR2_X1 U4045 ( .A1(n6633), .A2(n7053), .ZN(n4489) );
  OAI21_X2 U4046 ( .B1(n6652), .B2(n4495), .A(n3396), .ZN(n4496) );
  NOR2_X1 U4047 ( .A1(net218640), .A2(n4607), .ZN(n4475) );
  NOR2_X1 U4048 ( .A1(net216097), .A2(net218598), .ZN(n4474) );
  NOR2_X2 U4049 ( .A1(net212677), .A2(n4476), .ZN(n4480) );
  NOR2_X1 U4050 ( .A1(n3360), .A2(n4942), .ZN(n4198) );
  OAI21_X1 U4051 ( .B1(net215584), .B2(net218640), .A(net218610), .ZN(
        net217944) );
  NOR2_X2 U4052 ( .A1(net212677), .A2(n4004), .ZN(n4166) );
  NOR2_X2 U4053 ( .A1(b[9]), .A2(net218659), .ZN(n4004) );
  OAI21_X1 U4054 ( .B1(n4769), .B2(n4768), .A(n4767), .ZN(n4770) );
  NOR2_X1 U4055 ( .A1(n4777), .A2(n4942), .ZN(n4781) );
  NOR2_X1 U4056 ( .A1(net215210), .A2(net218598), .ZN(net217298) );
  NOR2_X1 U4057 ( .A1(net218640), .A2(net217299), .ZN(n4710) );
  NOR2_X2 U4058 ( .A1(net212677), .A2(n4711), .ZN(n4757) );
  NOR2_X2 U4059 ( .A1(b[10]), .A2(net218659), .ZN(n4711) );
  OAI21_X1 U4060 ( .B1(n7059), .B2(n5323), .A(n4857), .ZN(n4858) );
  AOI21_X2 U4061 ( .B1(n5174), .B2(n4865), .A(n4864), .ZN(n4866) );
  NOR2_X1 U4062 ( .A1(n4863), .A2(net218606), .ZN(n4864) );
  NOR2_X1 U4063 ( .A1(n5331), .A2(n3996), .ZN(n4869) );
  NOR2_X1 U4064 ( .A1(net218640), .A2(n4787), .ZN(n4789) );
  NOR2_X1 U4065 ( .A1(n6382), .A2(net218598), .ZN(n4788) );
  NOR2_X2 U4066 ( .A1(net212677), .A2(n4790), .ZN(n4847) );
  NOR2_X2 U4067 ( .A1(b[11]), .A2(net218659), .ZN(n4790) );
  NOR2_X1 U4068 ( .A1(net218640), .A2(n4875), .ZN(n4876) );
  OAI21_X1 U4069 ( .B1(n7078), .B2(n3338), .A(n3395), .ZN(n4955) );
  NOR2_X1 U4070 ( .A1(n7081), .A2(n7053), .ZN(n4944) );
  NOR2_X1 U4071 ( .A1(n4943), .A2(n4942), .ZN(n4945) );
  OAI21_X1 U4072 ( .B1(n7080), .B2(n6135), .A(n3392), .ZN(n4946) );
  NOR2_X2 U4073 ( .A1(net212677), .A2(n4878), .ZN(n4937) );
  NOR2_X2 U4074 ( .A1(b[12]), .A2(net218660), .ZN(n4878) );
  OAI21_X1 U4075 ( .B1(n3379), .B2(n5323), .A(n5048), .ZN(n5049) );
  NOR2_X1 U4076 ( .A1(n5058), .A2(n5332), .ZN(n5059) );
  AOI21_X2 U4077 ( .B1(n5174), .B2(n5054), .A(n5053), .ZN(n5055) );
  NOR2_X1 U4078 ( .A1(net216698), .A2(net218608), .ZN(n5053) );
  NOR2_X1 U4079 ( .A1(n5057), .A2(n3996), .ZN(n5061) );
  NOR2_X1 U4080 ( .A1(net216692), .A2(n5330), .ZN(n5060) );
  NOR2_X1 U4081 ( .A1(net213443), .A2(net218598), .ZN(net216855) );
  NOR2_X1 U4082 ( .A1(net218640), .A2(net216856), .ZN(n4961) );
  NOR2_X2 U4083 ( .A1(net212677), .A2(n4962), .ZN(n5036) );
  NOR2_X2 U4084 ( .A1(b[13]), .A2(net218660), .ZN(n4962) );
  OAI21_X1 U4085 ( .B1(n5169), .B2(n5323), .A(n5168), .ZN(n5170) );
  NOR2_X1 U4086 ( .A1(n5181), .A2(n5332), .ZN(n5182) );
  AOI21_X2 U4087 ( .B1(n5174), .B2(n7829), .A(n5173), .ZN(n5175) );
  NOR2_X1 U4088 ( .A1(n5172), .A2(net218606), .ZN(n5173) );
  NOR2_X2 U4089 ( .A1(n5179), .A2(n3996), .ZN(n5184) );
  NOR2_X1 U4090 ( .A1(n5180), .A2(n5330), .ZN(n5183) );
  NOR2_X1 U4091 ( .A1(n7246), .A2(net218598), .ZN(n5068) );
  NOR2_X1 U4092 ( .A1(net218640), .A2(n5067), .ZN(n5069) );
  NOR2_X2 U4093 ( .A1(net212677), .A2(n5070), .ZN(n5160) );
  NOR2_X2 U4094 ( .A1(b[14]), .A2(net218660), .ZN(n5070) );
  OAI21_X1 U4095 ( .B1(n7876), .B2(n5323), .A(n5322), .ZN(n5324) );
  NOR2_X1 U4096 ( .A1(net216306), .A2(n5332), .ZN(n5333) );
  NOR2_X1 U4097 ( .A1(n7041), .A2(n3996), .ZN(n5335) );
  NOR2_X1 U4098 ( .A1(n5331), .A2(n5330), .ZN(n5334) );
  NOR2_X1 U4099 ( .A1(n7589), .A2(net218600), .ZN(n5191) );
  NOR2_X1 U4100 ( .A1(net218640), .A2(n5190), .ZN(n5192) );
  NOR2_X2 U4101 ( .A1(net212677), .A2(n5194), .ZN(n5309) );
  NOR2_X2 U4102 ( .A1(b[15]), .A2(net218660), .ZN(n5194) );
  NOR2_X1 U4103 ( .A1(n6144), .A2(net218640), .ZN(n6146) );
  NOR2_X1 U4104 ( .A1(net214758), .A2(net218608), .ZN(n6145) );
  NOR2_X1 U4105 ( .A1(n6277), .A2(n6984), .ZN(n6281) );
  NOR2_X1 U4106 ( .A1(n6279), .A2(n6983), .ZN(n6280) );
  OAI21_X1 U4107 ( .B1(n6638), .B2(n7058), .A(n3385), .ZN(n6640) );
  NOR2_X2 U4108 ( .A1(n6635), .A2(n6634), .ZN(n6638) );
  OAI21_X1 U4109 ( .B1(n6633), .B2(n3993), .A(n3391), .ZN(n6634) );
  OAI21_X1 U4110 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(n6654) );
  NOR2_X1 U4111 ( .A1(net214219), .A2(net218610), .ZN(n6655) );
  NOR2_X2 U4112 ( .A1(n5456), .A2(n3372), .ZN(n5458) );
  NOR2_X1 U4113 ( .A1(n7080), .A2(n6983), .ZN(n6628) );
  NOR2_X1 U4114 ( .A1(n7381), .A2(n7828), .ZN(n7391) );
  NOR2_X2 U4115 ( .A1(n7389), .A2(n7388), .ZN(n7390) );
  NOR2_X2 U4116 ( .A1(n7232), .A2(n7231), .ZN(n7394) );
  NOR2_X1 U4117 ( .A1(n7230), .A2(net218640), .ZN(n7231) );
  AOI21_X1 U4118 ( .B1(n7229), .B2(n7228), .A(n7878), .ZN(n7232) );
  OAI21_X1 U4119 ( .B1(n7220), .B2(n3390), .A(n7866), .ZN(n7229) );
  INV_X4 U4120 ( .A(net212097), .ZN(net223578) );
  OAI21_X1 U4121 ( .B1(b[31]), .B2(net218660), .A(net212094), .ZN(net212097)
         );
  AOI21_X1 U4122 ( .B1(net212677), .B2(n4274), .A(n4262), .ZN(n4291) );
  AOI211_X2 U4123 ( .C1(n5452), .C2(n5588), .A(n3386), .B(n6639), .ZN(n5466)
         );
  AOI222_X1 U4124 ( .A1(n6851), .A2(n6850), .B1(n7031), .B2(n5595), .C1(n7033), 
        .C2(n6123), .ZN(n5612) );
  AOI222_X1 U4125 ( .A1(n6851), .A2(n6982), .B1(n7031), .B2(n5739), .C1(n7033), 
        .C2(n6278), .ZN(n5755) );
  AOI222_X1 U4126 ( .A1(n6851), .A2(net213359), .B1(n7031), .B2(n6451), .C1(
        n7033), .C2(net214477), .ZN(n5884) );
  NAND3_X2 U4127 ( .A1(n6011), .A2(n6010), .A3(n6009), .ZN(result[20]) );
  AOI211_X2 U4128 ( .C1(b[20]), .C2(n5991), .A(n5990), .B(n5989), .ZN(n6011)
         );
  NAND3_X2 U4129 ( .A1(n6130), .A2(n6129), .A3(n6128), .ZN(result[21]) );
  NAND3_X2 U4130 ( .A1(n6482), .A2(n6481), .A3(n6480), .ZN(result[23]) );
  AOI211_X2 U4131 ( .C1(b[23]), .C2(n6479), .A(n6478), .B(n6477), .ZN(n6480)
         );
  AOI222_X1 U4132 ( .A1(n6851), .A2(n7222), .B1(n7031), .B2(n6850), .C1(n7033), 
        .C2(n6849), .ZN(n6866) );
  NOR3_X2 U4133 ( .A1(n6988), .A2(n6987), .A3(n6986), .ZN(n7008) );
  AOI211_X2 U4134 ( .C1(n7045), .C2(n7044), .A(n7043), .B(n7042), .ZN(n7064)
         );
  AOI21_X1 U4135 ( .B1(n7099), .B2(n7098), .A(net213275), .ZN(n7212) );
  AOI21_X1 U4136 ( .B1(n7091), .B2(n7821), .A(n7090), .ZN(n7214) );
  NOR2_X1 U4137 ( .A1(n7892), .A2(n7891), .ZN(n7894) );
  INV_X8 U4138 ( .A(n3365), .ZN(n3990) );
  INV_X16 U4139 ( .A(a[8]), .ZN(net218434) );
  INV_X16 U4140 ( .A(a[9]), .ZN(net218428) );
  INV_X16 U4141 ( .A(a[11]), .ZN(net218414) );
  INV_X16 U4142 ( .A(a[15]), .ZN(n3487) );
  INV_X4 U4143 ( .A(sel), .ZN(n4001) );
  INV_X16 U4144 ( .A(b[6]), .ZN(n3485) );
  AND2_X4 U4145 ( .A1(b[5]), .A2(a[15]), .ZN(n3303) );
  INV_X16 U4146 ( .A(b[11]), .ZN(n3486) );
  AND2_X4 U4147 ( .A1(a[22]), .A2(b[6]), .ZN(n3304) );
  INV_X16 U4148 ( .A(b[13]), .ZN(net218502) );
  INV_X16 U4149 ( .A(a[12]), .ZN(net218406) );
  INV_X16 U4150 ( .A(a[13]), .ZN(net218400) );
  INV_X16 U4151 ( .A(a[14]), .ZN(net218392) );
  INV_X8 U4152 ( .A(a[1]), .ZN(net218484) );
  INV_X4 U4153 ( .A(net218484), .ZN(net218480) );
  AND2_X2 U4154 ( .A1(net218550), .A2(a[0]), .ZN(n3305) );
  OR2_X2 U4155 ( .A1(result[28]), .A2(n3349), .ZN(n3306) );
  INV_X16 U4156 ( .A(a[10]), .ZN(net218420) );
  AND2_X4 U4157 ( .A1(b[5]), .A2(a[12]), .ZN(n3307) );
  AND2_X2 U4158 ( .A1(b[5]), .A2(a[8]), .ZN(n3308) );
  AND2_X4 U4159 ( .A1(b[4]), .A2(a[15]), .ZN(n3309) );
  AND2_X4 U4160 ( .A1(b[4]), .A2(a[16]), .ZN(n3310) );
  AND2_X4 U4161 ( .A1(a[13]), .A2(b[4]), .ZN(n3311) );
  AND2_X4 U4162 ( .A1(b[5]), .A2(a[9]), .ZN(n3312) );
  AND2_X4 U4163 ( .A1(b[7]), .A2(a[3]), .ZN(n3313) );
  AND2_X4 U4164 ( .A1(b[4]), .A2(a[11]), .ZN(n3314) );
  AND2_X4 U4165 ( .A1(b[5]), .A2(a[11]), .ZN(n3315) );
  AND2_X4 U4166 ( .A1(b[7]), .A2(net218480), .ZN(n3316) );
  AND2_X2 U4167 ( .A1(b[4]), .A2(a[17]), .ZN(n3317) );
  OR2_X4 U4168 ( .A1(result[24]), .A2(n3346), .ZN(n3318) );
  OR2_X2 U4169 ( .A1(result[22]), .A2(n3348), .ZN(n3319) );
  OR2_X2 U4170 ( .A1(result[26]), .A2(n3345), .ZN(n3320) );
  AND2_X4 U4171 ( .A1(a[13]), .A2(b[6]), .ZN(n3321) );
  AND2_X4 U4172 ( .A1(b[8]), .A2(a[9]), .ZN(n3322) );
  AND2_X4 U4173 ( .A1(a[22]), .A2(b[7]), .ZN(n3323) );
  AND2_X4 U4174 ( .A1(a[24]), .A2(b[5]), .ZN(n3324) );
  OR2_X2 U4175 ( .A1(result[14]), .A2(n3359), .ZN(n3325) );
  OR2_X2 U4176 ( .A1(result[19]), .A2(n3352), .ZN(n3326) );
  AND2_X4 U4177 ( .A1(b[17]), .A2(net219055), .ZN(n3327) );
  AND2_X4 U4178 ( .A1(a[16]), .A2(b[12]), .ZN(n3328) );
  OR2_X2 U4179 ( .A1(b[4]), .A2(net219055), .ZN(n3329) );
  OR2_X2 U4180 ( .A1(result[6]), .A2(n3388), .ZN(n3330) );
  AND2_X4 U4181 ( .A1(a[2]), .A2(b[27]), .ZN(n3331) );
  INV_X8 U4182 ( .A(net211994), .ZN(net218639) );
  AND2_X2 U4183 ( .A1(n3998), .A2(a[24]), .ZN(n3332) );
  XOR2_X2 U4184 ( .A(n5871), .B(net215709), .Z(n3334) );
  XOR2_X2 U4185 ( .A(n6105), .B(net215252), .Z(n3335) );
  XOR2_X2 U4186 ( .A(n6852), .B(net214219), .Z(n3336) );
  XOR2_X2 U4187 ( .A(n7047), .B(n6999), .Z(n3337) );
  OR2_X4 U4188 ( .A1(net218544), .A2(n5323), .ZN(n3338) );
  INV_X4 U4189 ( .A(n4001), .ZN(n4002) );
  INV_X4 U4190 ( .A(n3888), .ZN(n3978) );
  INV_X4 U4191 ( .A(net217295), .ZN(net217233) );
  AND2_X2 U4192 ( .A1(n7627), .A2(n7459), .ZN(n3340) );
  INV_X4 U4193 ( .A(net215057), .ZN(n3700) );
  OR2_X2 U4194 ( .A1(net217135), .A2(net217136), .ZN(n3341) );
  INV_X4 U4195 ( .A(n5585), .ZN(n5586) );
  AND2_X2 U4196 ( .A1(n3299), .A2(net216985), .ZN(n3342) );
  AND2_X2 U4197 ( .A1(a[3]), .A2(a[4]), .ZN(n3343) );
  INV_X16 U4198 ( .A(a[2]), .ZN(net218476) );
  XOR2_X1 U4199 ( .A(n7524), .B(n7758), .Z(n3344) );
  OR2_X2 U4200 ( .A1(result[25]), .A2(n3318), .ZN(n3345) );
  OR2_X2 U4201 ( .A1(result[23]), .A2(n3319), .ZN(n3346) );
  OR2_X2 U4202 ( .A1(result[20]), .A2(n3326), .ZN(n3347) );
  OR2_X2 U4203 ( .A1(result[21]), .A2(n3347), .ZN(n3348) );
  INV_X4 U4204 ( .A(net217083), .ZN(net219116) );
  OR2_X2 U4205 ( .A1(result[27]), .A2(n3320), .ZN(n3349) );
  INV_X4 U4206 ( .A(n5204), .ZN(n3814) );
  INV_X2 U4207 ( .A(n5298), .ZN(n5552) );
  AND2_X2 U4208 ( .A1(b[9]), .A2(a[2]), .ZN(n3350) );
  OR2_X2 U4209 ( .A1(result[15]), .A2(n3325), .ZN(n3351) );
  OR2_X2 U4210 ( .A1(result[18]), .A2(n3468), .ZN(n3352) );
  INV_X4 U4211 ( .A(n6382), .ZN(n3590) );
  INV_X4 U4212 ( .A(net216097), .ZN(net219220) );
  AND2_X4 U4213 ( .A1(b[15]), .A2(a[9]), .ZN(n3353) );
  XOR2_X2 U4214 ( .A(net217984), .B(a[6]), .Z(n3354) );
  AND3_X4 U4215 ( .A1(n7885), .A2(n7884), .A3(n7883), .ZN(n3355) );
  OR2_X2 U4216 ( .A1(result[7]), .A2(n3330), .ZN(n3356) );
  OR2_X2 U4217 ( .A1(result[9]), .A2(n7839), .ZN(n3357) );
  OR2_X2 U4218 ( .A1(result[10]), .A2(n3357), .ZN(n3358) );
  OR2_X2 U4219 ( .A1(result[13]), .A2(n7887), .ZN(n3359) );
  INV_X4 U4220 ( .A(net214293), .ZN(n3602) );
  INV_X4 U4221 ( .A(n3880), .ZN(n3988) );
  INV_X8 U4222 ( .A(n7869), .ZN(n7807) );
  AND4_X4 U4223 ( .A1(net216710), .A2(net216328), .A3(net217942), .A4(
        net217027), .ZN(n3360) );
  AND2_X4 U4224 ( .A1(b[24]), .A2(a[3]), .ZN(n3361) );
  AND2_X2 U4225 ( .A1(a[11]), .A2(b[19]), .ZN(n3362) );
  AND2_X4 U4226 ( .A1(b[27]), .A2(net218480), .ZN(n3363) );
  AND2_X4 U4227 ( .A1(n6003), .A2(n6002), .ZN(n3364) );
  AND2_X4 U4228 ( .A1(n3158), .A2(n4003), .ZN(n3365) );
  AND2_X2 U4229 ( .A1(n3997), .A2(a[14]), .ZN(n3366) );
  AND2_X4 U4230 ( .A1(n3997), .A2(a[18]), .ZN(n3367) );
  AND2_X4 U4231 ( .A1(n3997), .A2(a[22]), .ZN(n3368) );
  AND2_X4 U4232 ( .A1(n4345), .A2(n4416), .ZN(n3369) );
  AND2_X4 U4233 ( .A1(b[25]), .A2(a[1]), .ZN(n3370) );
  AND2_X2 U4234 ( .A1(n3997), .A2(a[26]), .ZN(n3371) );
  AND2_X2 U4235 ( .A1(n3998), .A2(a[16]), .ZN(n3372) );
  AND2_X2 U4236 ( .A1(n3998), .A2(a[20]), .ZN(n3373) );
  INV_X16 U4237 ( .A(net211950), .ZN(net218614) );
  AND2_X2 U4238 ( .A1(n3998), .A2(a[8]), .ZN(n3374) );
  AND2_X2 U4239 ( .A1(n3998), .A2(a[12]), .ZN(n3375) );
  AND2_X4 U4240 ( .A1(b[21]), .A2(a[2]), .ZN(n3376) );
  OAI21_X2 U4241 ( .B1(net218558), .B2(n4700), .A(n4267), .ZN(n6100) );
  AND2_X4 U4242 ( .A1(n7807), .A2(n4235), .ZN(n3377) );
  INV_X1 U4243 ( .A(n6982), .ZN(n6277) );
  XOR2_X2 U4244 ( .A(a[18]), .B(b[18]), .Z(n3378) );
  AND2_X4 U4245 ( .A1(n5047), .A2(n5046), .ZN(n3379) );
  OR2_X4 U4246 ( .A1(net218534), .A2(n7035), .ZN(n3380) );
  OR2_X4 U4247 ( .A1(net218534), .A2(n7058), .ZN(n3381) );
  AND2_X2 U4248 ( .A1(n5736), .A2(n6272), .ZN(n3382) );
  INV_X16 U4249 ( .A(net212100), .ZN(net218658) );
  OR2_X2 U4250 ( .A1(net218534), .A2(n5323), .ZN(n3383) );
  AND2_X2 U4251 ( .A1(n5736), .A2(n6100), .ZN(n3384) );
  OR2_X4 U4252 ( .A1(n6637), .A2(n6636), .ZN(n3385) );
  AND2_X2 U4253 ( .A1(n5736), .A2(n5451), .ZN(n3386) );
  OR2_X2 U4254 ( .A1(result[4]), .A2(n7836), .ZN(n3387) );
  OR2_X2 U4255 ( .A1(result[5]), .A2(n3387), .ZN(n3388) );
  AND2_X2 U4256 ( .A1(n7031), .A2(net213359), .ZN(n3389) );
  OR2_X4 U4257 ( .A1(n7219), .A2(n7218), .ZN(n3390) );
  OR2_X4 U4258 ( .A1(n3995), .A2(n6632), .ZN(n3391) );
  OR2_X4 U4259 ( .A1(net214022), .A2(net218598), .ZN(n3392) );
  OR2_X2 U4260 ( .A1(net218534), .A2(n4860), .ZN(n3393) );
  OR2_X4 U4261 ( .A1(net217244), .A2(net218598), .ZN(n3394) );
  OR2_X4 U4262 ( .A1(n4951), .A2(net218606), .ZN(n3395) );
  OR2_X4 U4263 ( .A1(n4494), .A2(net218606), .ZN(n3396) );
  INV_X16 U4264 ( .A(net211949), .ZN(net218604) );
  OR2_X4 U4265 ( .A1(net215799), .A2(net218600), .ZN(n3397) );
  OR2_X4 U4266 ( .A1(net215709), .A2(net218600), .ZN(n3398) );
  OR2_X4 U4267 ( .A1(net215709), .A2(net218608), .ZN(n3399) );
  OR2_X4 U4268 ( .A1(net216124), .A2(net218600), .ZN(n3400) );
  OR2_X4 U4269 ( .A1(net216124), .A2(net218608), .ZN(n3401) );
  OR2_X4 U4270 ( .A1(net215252), .A2(net218608), .ZN(n3402) );
  OR2_X4 U4271 ( .A1(net215499), .A2(net218600), .ZN(n3403) );
  OR2_X4 U4272 ( .A1(net215499), .A2(net218608), .ZN(n3404) );
  OR2_X4 U4273 ( .A1(net213919), .A2(net218600), .ZN(n3405) );
  OR2_X4 U4274 ( .A1(n7054), .A2(net218600), .ZN(n3406) );
  OR2_X4 U4275 ( .A1(n6999), .A2(net218600), .ZN(n3407) );
  OR2_X4 U4276 ( .A1(net217796), .A2(net218606), .ZN(n3408) );
  OR2_X4 U4277 ( .A1(n5328), .A2(net218608), .ZN(n3409) );
  OR2_X4 U4278 ( .A1(net217169), .A2(net218606), .ZN(n3410) );
  INV_X16 U4279 ( .A(n3992), .ZN(n3993) );
  INV_X4 U4280 ( .A(n7870), .ZN(n3992) );
  OR2_X4 U4281 ( .A1(net218484), .A2(net218598), .ZN(n3411) );
  OR2_X4 U4282 ( .A1(net218378), .A2(net218600), .ZN(n3412) );
  OR2_X4 U4283 ( .A1(net215252), .A2(net218600), .ZN(n3413) );
  OR2_X4 U4284 ( .A1(net214219), .A2(net218600), .ZN(n3414) );
  INV_X4 U4285 ( .A(n4001), .ZN(n4000) );
  OAI21_X2 U4286 ( .B1(n5614), .B2(n5615), .A(n5892), .ZN(n5710) );
  OAI21_X2 U4287 ( .B1(net214427), .B2(net214428), .A(net214429), .ZN(n6511)
         );
  NAND2_X2 U4288 ( .A1(n3843), .A2(n3840), .ZN(n3848) );
  INV_X8 U4289 ( .A(net214025), .ZN(net213870) );
  XNOR2_X2 U4290 ( .A(n6824), .B(n6823), .ZN(n3924) );
  INV_X2 U4291 ( .A(n5212), .ZN(n3415) );
  INV_X4 U4292 ( .A(n3415), .ZN(n3416) );
  XNOR2_X2 U4293 ( .A(n5844), .B(n5849), .ZN(n3417) );
  AOI21_X4 U4294 ( .B1(net214877), .B2(net214878), .A(net214879), .ZN(
        net215122) );
  NAND2_X2 U4295 ( .A1(n7010), .A2(n7104), .ZN(n6973) );
  NAND2_X4 U4296 ( .A1(n6971), .A2(n3370), .ZN(n7104) );
  NAND2_X4 U4297 ( .A1(n3582), .A2(n3583), .ZN(net215061) );
  XNOR2_X2 U4298 ( .A(n6781), .B(net214033), .ZN(n3418) );
  NAND2_X2 U4299 ( .A1(n6197), .A2(n6196), .ZN(n6519) );
  INV_X2 U4300 ( .A(n6196), .ZN(n6194) );
  NAND2_X2 U4301 ( .A1(n6171), .A2(n6170), .ZN(n6334) );
  NAND2_X4 U4302 ( .A1(n6366), .A2(n6365), .ZN(n6726) );
  INV_X2 U4303 ( .A(n4880), .ZN(n3922) );
  INV_X8 U4304 ( .A(net215331), .ZN(net214963) );
  NAND2_X2 U4305 ( .A1(net213227), .A2(net213225), .ZN(net213414) );
  XNOR2_X2 U4306 ( .A(n5426), .B(n3886), .ZN(n5427) );
  NAND2_X4 U4307 ( .A1(net213396), .A2(net220449), .ZN(net212942) );
  XNOR2_X2 U4308 ( .A(n6788), .B(net219938), .ZN(n6789) );
  NAND2_X4 U4309 ( .A1(n6956), .A2(n3195), .ZN(net213680) );
  INV_X4 U4310 ( .A(net217790), .ZN(net217857) );
  NAND2_X2 U4311 ( .A1(net217243), .A2(net216946), .ZN(net218066) );
  OAI21_X2 U4312 ( .B1(n4016), .B2(n3763), .A(n4015), .ZN(n4012) );
  OAI21_X4 U4313 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(n4109) );
  XNOR2_X2 U4314 ( .A(n5143), .B(n5142), .ZN(n3419) );
  NAND2_X2 U4315 ( .A1(n5904), .A2(n5626), .ZN(n5549) );
  INV_X2 U4316 ( .A(net214570), .ZN(net214830) );
  NAND2_X4 U4317 ( .A1(net214571), .A2(net220181), .ZN(n6244) );
  NOR2_X2 U4318 ( .A1(n3689), .A2(n3690), .ZN(net216573) );
  INV_X4 U4319 ( .A(n6012), .ZN(n5888) );
  INV_X2 U4320 ( .A(net218109), .ZN(n3420) );
  INV_X2 U4321 ( .A(n6880), .ZN(n3421) );
  INV_X2 U4322 ( .A(n6878), .ZN(n6880) );
  INV_X4 U4323 ( .A(n5231), .ZN(n5234) );
  OAI211_X4 U4324 ( .C1(n5353), .C2(net216277), .A(n5352), .B(net216279), .ZN(
        n5477) );
  NAND2_X2 U4325 ( .A1(n5351), .A2(net216284), .ZN(n5220) );
  NAND2_X4 U4326 ( .A1(n5475), .A2(n5474), .ZN(n5639) );
  NAND3_X2 U4327 ( .A1(a[0]), .A2(b[11]), .A3(n4934), .ZN(n3422) );
  NAND2_X4 U4328 ( .A1(net212951), .A2(net212655), .ZN(n3423) );
  NAND2_X4 U4329 ( .A1(n7024), .A2(n3361), .ZN(net212655) );
  OAI21_X4 U4330 ( .B1(n4970), .B2(n4969), .A(n4968), .ZN(n5207) );
  NAND2_X2 U4331 ( .A1(n5536), .A2(n5535), .ZN(net215674) );
  NAND2_X2 U4332 ( .A1(n5978), .A2(n5979), .ZN(net214983) );
  XNOR2_X2 U4333 ( .A(net214792), .B(net214793), .ZN(n3424) );
  NAND2_X2 U4334 ( .A1(n7024), .A2(n3361), .ZN(n3425) );
  XNOR2_X2 U4335 ( .A(n6418), .B(n6417), .ZN(n3426) );
  NAND2_X2 U4336 ( .A1(n6673), .A2(n6873), .ZN(n6874) );
  XNOR2_X2 U4337 ( .A(net215571), .B(n5823), .ZN(n3427) );
  AOI21_X4 U4338 ( .B1(net215775), .B2(n3764), .A(n3787), .ZN(n5823) );
  AOI21_X2 U4339 ( .B1(b[28]), .B2(n7210), .A(n7209), .ZN(n7211) );
  INV_X2 U4340 ( .A(net212404), .ZN(n3428) );
  INV_X4 U4341 ( .A(n3428), .ZN(n3429) );
  NAND2_X4 U4342 ( .A1(net218146), .A2(net218147), .ZN(net217292) );
  NAND3_X2 U4343 ( .A1(n7393), .A2(n7392), .A3(n7394), .ZN(result[29]) );
  NAND4_X2 U4344 ( .A1(net211939), .A2(n7893), .A3(net223581), .A4(n7894), 
        .ZN(result[30]) );
  NAND2_X2 U4345 ( .A1(net213423), .A2(net213422), .ZN(net213221) );
  OAI21_X4 U4346 ( .B1(net213219), .B2(net213220), .A(net213221), .ZN(
        net212916) );
  INV_X4 U4347 ( .A(net213421), .ZN(net213423) );
  NAND2_X4 U4348 ( .A1(net213420), .A2(net213421), .ZN(net213223) );
  INV_X4 U4349 ( .A(net213422), .ZN(net213420) );
  NAND2_X4 U4350 ( .A1(net212643), .A2(net212731), .ZN(net213017) );
  XNOR2_X2 U4351 ( .A(net213017), .B(net213018), .ZN(net213013) );
  NAND2_X4 U4352 ( .A1(net213028), .A2(net213027), .ZN(net212643) );
  INV_X4 U4353 ( .A(net213026), .ZN(net213028) );
  NAND2_X1 U4354 ( .A1(net213027), .A2(net213028), .ZN(net219746) );
  XNOR2_X2 U4355 ( .A(net213029), .B(net213030), .ZN(net213026) );
  NAND2_X4 U4356 ( .A1(net219933), .A2(net213025), .ZN(net212731) );
  INV_X1 U4357 ( .A(net212731), .ZN(net212644) );
  INV_X4 U4358 ( .A(net213027), .ZN(net213025) );
  XNOR2_X2 U4359 ( .A(net213029), .B(net213030), .ZN(net219933) );
  NAND2_X2 U4360 ( .A1(b[22]), .A2(a[6]), .ZN(net213027) );
  NAND2_X4 U4361 ( .A1(net212941), .A2(net219504), .ZN(net213030) );
  INV_X2 U4362 ( .A(net219503), .ZN(net219504) );
  INV_X2 U4363 ( .A(net212942), .ZN(net219503) );
  OAI21_X2 U4364 ( .B1(net213031), .B2(n3208), .A(net213033), .ZN(net212941)
         );
  NOR2_X4 U4365 ( .A1(net213031), .A2(n3208), .ZN(net213391) );
  INV_X4 U4366 ( .A(net213603), .ZN(net213600) );
  XOR2_X1 U4367 ( .A(net213700), .B(net213701), .Z(n3431) );
  NAND2_X4 U4368 ( .A1(net219693), .A2(net213036), .ZN(net212938) );
  INV_X4 U4369 ( .A(net212935), .ZN(net212933) );
  OAI21_X4 U4370 ( .B1(net212933), .B2(net212932), .A(net212934), .ZN(
        net212470) );
  NAND2_X4 U4371 ( .A1(net213035), .A2(net213034), .ZN(net212940) );
  NAND2_X4 U4372 ( .A1(n3432), .A2(net212422), .ZN(net212424) );
  XNOR2_X2 U4373 ( .A(net212424), .B(n3331), .ZN(net212423) );
  NAND2_X4 U4374 ( .A1(net212710), .A2(net212709), .ZN(n3432) );
  INV_X4 U4375 ( .A(net219333), .ZN(net212710) );
  NAND2_X2 U4376 ( .A1(net212709), .A2(net212710), .ZN(net220061) );
  XNOR2_X2 U4377 ( .A(net224024), .B(net212711), .ZN(net219333) );
  INV_X4 U4378 ( .A(net219421), .ZN(net212445) );
  NAND2_X4 U4379 ( .A1(net212445), .A2(net212439), .ZN(net224024) );
  NAND2_X4 U4380 ( .A1(net212708), .A2(net212707), .ZN(net212422) );
  NAND2_X4 U4381 ( .A1(net212422), .A2(net220061), .ZN(net212420) );
  BUF_X8 U4382 ( .A(net212422), .Z(net220011) );
  INV_X4 U4383 ( .A(net212709), .ZN(net212707) );
  XNOR2_X2 U4384 ( .A(net224024), .B(net212711), .ZN(net212708) );
  NAND2_X2 U4385 ( .A1(a[3]), .A2(b[26]), .ZN(net212709) );
  NAND2_X4 U4386 ( .A1(net212442), .A2(net219464), .ZN(net212711) );
  INV_X4 U4387 ( .A(net219463), .ZN(net219464) );
  AOI21_X1 U4388 ( .B1(net212442), .B2(net219464), .A(net219421), .ZN(
        net212437) );
  INV_X2 U4389 ( .A(net212443), .ZN(net219463) );
  NAND2_X4 U4390 ( .A1(net212440), .A2(net212441), .ZN(net212439) );
  CLKBUF_X3 U4391 ( .A(net212439), .Z(net223689) );
  XNOR2_X2 U4392 ( .A(net212714), .B(net212713), .ZN(net212440) );
  XNOR2_X2 U4393 ( .A(net219422), .B(net212717), .ZN(net219421) );
  NAND3_X2 U4394 ( .A1(net212648), .A2(net212647), .A3(net212718), .ZN(
        net212717) );
  INV_X4 U4395 ( .A(net212441), .ZN(net212718) );
  AND2_X2 U4396 ( .A1(net212715), .A2(net212718), .ZN(net219422) );
  NAND2_X2 U4397 ( .A1(net212954), .A2(net212443), .ZN(net213000) );
  NOR2_X1 U4398 ( .A1(net219357), .A2(net212441), .ZN(net212438) );
  XNOR2_X1 U4399 ( .A(net212714), .B(net212713), .ZN(net219357) );
  NAND2_X4 U4400 ( .A1(net212648), .A2(net212647), .ZN(net212714) );
  NAND2_X4 U4401 ( .A1(net216802), .A2(net216803), .ZN(net216801) );
  INV_X4 U4402 ( .A(net216801), .ZN(net216798) );
  NAND2_X4 U4403 ( .A1(net217124), .A2(net217125), .ZN(net216802) );
  OAI21_X1 U4404 ( .B1(net217125), .B2(net217124), .A(net216802), .ZN(
        net217121) );
  NAND2_X2 U4405 ( .A1(net216803), .A2(net216802), .ZN(net216961) );
  INV_X4 U4406 ( .A(net217126), .ZN(net217125) );
  NAND2_X2 U4407 ( .A1(net216966), .A2(net216967), .ZN(net216803) );
  INV_X4 U4408 ( .A(net216968), .ZN(net216967) );
  INV_X2 U4409 ( .A(net216517), .ZN(net216966) );
  XNOR2_X2 U4410 ( .A(net216968), .B(net216517), .ZN(net217126) );
  NAND2_X4 U4411 ( .A1(net216448), .A2(net216449), .ZN(net216447) );
  INV_X4 U4412 ( .A(net216447), .ZN(net216444) );
  NAND2_X4 U4413 ( .A1(n3433), .A2(net216628), .ZN(net216448) );
  NAND2_X2 U4414 ( .A1(net216449), .A2(net216448), .ZN(net216623) );
  INV_X4 U4415 ( .A(net216797), .ZN(net216628) );
  OAI22_X2 U4416 ( .A1(net216628), .A2(net219485), .B1(net216796), .B2(
        net216797), .ZN(net216794) );
  OAI21_X4 U4417 ( .B1(net216798), .B2(net216799), .A(net216800), .ZN(n3433)
         );
  OAI21_X2 U4418 ( .B1(net216798), .B2(net216799), .A(net216800), .ZN(
        net219485) );
  NAND2_X2 U4419 ( .A1(net216630), .A2(net216631), .ZN(net216449) );
  INV_X4 U4420 ( .A(net216632), .ZN(net216631) );
  INV_X4 U4421 ( .A(net216117), .ZN(net216630) );
  XNOR2_X2 U4422 ( .A(net216961), .B(net216799), .ZN(net216958) );
  NAND2_X2 U4423 ( .A1(net216962), .A2(net216800), .ZN(net216799) );
  XNOR2_X2 U4424 ( .A(net216632), .B(net216117), .ZN(net216797) );
  NAND2_X4 U4425 ( .A1(net216074), .A2(net216075), .ZN(net216073) );
  INV_X4 U4426 ( .A(net216073), .ZN(net216070) );
  NAND2_X4 U4427 ( .A1(net216442), .A2(net216441), .ZN(net216074) );
  OAI21_X2 U4428 ( .B1(net216442), .B2(net216441), .A(net216074), .ZN(
        net216439) );
  NAND2_X4 U4429 ( .A1(net216074), .A2(net216075), .ZN(net216252) );
  INV_X4 U4430 ( .A(net216443), .ZN(net216442) );
  NAND2_X2 U4431 ( .A1(net216257), .A2(net216258), .ZN(net216075) );
  INV_X4 U4432 ( .A(net216259), .ZN(net216258) );
  INV_X4 U4433 ( .A(net215701), .ZN(net216257) );
  XNOR2_X2 U4434 ( .A(net216259), .B(net215701), .ZN(net216443) );
  NAND2_X4 U4435 ( .A1(net212924), .A2(net212926), .ZN(net213048) );
  XNOR2_X2 U4436 ( .A(net213048), .B(n3161), .ZN(net213046) );
  OAI21_X4 U4437 ( .B1(net212922), .B2(net212923), .A(net212924), .ZN(
        net212485) );
  XNOR2_X2 U4438 ( .A(net213053), .B(net213054), .ZN(net220068) );
  INV_X4 U4439 ( .A(net212919), .ZN(net213053) );
  XNOR2_X2 U4440 ( .A(net213053), .B(net213054), .ZN(n3434) );
  INV_X4 U4441 ( .A(net213050), .ZN(net213052) );
  NAND2_X4 U4442 ( .A1(net213049), .A2(net213050), .ZN(net212926) );
  INV_X4 U4443 ( .A(n3434), .ZN(net213049) );
  OAI21_X2 U4444 ( .B1(net212918), .B2(net212919), .A(net212920), .ZN(
        net212495) );
  NAND2_X4 U4445 ( .A1(net212929), .A2(net212931), .ZN(net213043) );
  XNOR2_X2 U4446 ( .A(net212930), .B(net213043), .ZN(net213041) );
  NAND2_X2 U4447 ( .A1(net213046), .A2(net213047), .ZN(net212929) );
  INV_X4 U4448 ( .A(net213045), .ZN(net213047) );
  NAND2_X4 U4449 ( .A1(net213044), .A2(net213045), .ZN(net212931) );
  INV_X2 U4450 ( .A(net212931), .ZN(net212927) );
  INV_X4 U4451 ( .A(net213046), .ZN(net213044) );
  NAND2_X4 U4452 ( .A1(net213216), .A2(net213218), .ZN(net213424) );
  XNOR2_X2 U4453 ( .A(net213217), .B(net213424), .ZN(net213422) );
  NAND2_X4 U4454 ( .A1(net213427), .A2(net213428), .ZN(net213216) );
  OAI21_X4 U4455 ( .B1(net213214), .B2(net213215), .A(net213216), .ZN(
        net212911) );
  INV_X4 U4456 ( .A(net213426), .ZN(net213428) );
  XNOR2_X2 U4457 ( .A(net213212), .B(net213429), .ZN(net213427) );
  NAND2_X4 U4458 ( .A1(net224071), .A2(net213426), .ZN(net213218) );
  INV_X1 U4459 ( .A(net213218), .ZN(net213214) );
  XNOR2_X2 U4460 ( .A(net213429), .B(net213210), .ZN(net224071) );
  OAI21_X4 U4461 ( .B1(net213209), .B2(net213210), .A(net213211), .ZN(
        net213070) );
  NAND3_X1 U4462 ( .A1(net212650), .A2(net212649), .A3(net212648), .ZN(
        net212646) );
  INV_X1 U4463 ( .A(net212647), .ZN(net219678) );
  NAND2_X2 U4464 ( .A1(net212715), .A2(net212652), .ZN(net212713) );
  NAND2_X4 U4465 ( .A1(net213194), .A2(net212899), .ZN(net213455) );
  NAND2_X4 U4466 ( .A1(net213459), .A2(net213458), .ZN(net213194) );
  OAI21_X4 U4467 ( .B1(net213192), .B2(net213193), .A(net213194), .ZN(
        net212900) );
  INV_X4 U4468 ( .A(net213457), .ZN(net213459) );
  NAND2_X2 U4469 ( .A1(net213457), .A2(net213456), .ZN(net212899) );
  CLKBUF_X2 U4470 ( .A(net212899), .Z(net220199) );
  INV_X4 U4471 ( .A(net213458), .ZN(net213456) );
  INV_X4 U4472 ( .A(net213036), .ZN(net213034) );
  XNOR2_X2 U4473 ( .A(net213038), .B(net212935), .ZN(net213035) );
  NAND2_X4 U4474 ( .A1(net213033), .A2(net212942), .ZN(net213392) );
  NOR2_X4 U4475 ( .A1(n3436), .A2(net213174), .ZN(n3435) );
  XNOR2_X2 U4476 ( .A(n3435), .B(net213472), .ZN(net213469) );
  INV_X4 U4477 ( .A(net213475), .ZN(net213174) );
  OAI21_X1 U4478 ( .B1(net213174), .B2(net213472), .A(net213176), .ZN(
        net212883) );
  NAND2_X2 U4479 ( .A1(net219974), .A2(net213477), .ZN(net213475) );
  INV_X4 U4480 ( .A(net213176), .ZN(n3436) );
  XNOR2_X2 U4481 ( .A(net213170), .B(net213480), .ZN(net219974) );
  INV_X4 U4482 ( .A(net219974), .ZN(net213478) );
  NAND2_X2 U4483 ( .A1(net213171), .A2(net213173), .ZN(net213480) );
  INV_X4 U4484 ( .A(net213172), .ZN(net213170) );
  OAI21_X4 U4485 ( .B1(net213169), .B2(net213170), .A(net213171), .ZN(
        net212826) );
  OAI21_X4 U4486 ( .B1(n3437), .B2(n3438), .A(net213537), .ZN(net213172) );
  INV_X4 U4487 ( .A(net213538), .ZN(n3438) );
  INV_X4 U4488 ( .A(net213539), .ZN(n3437) );
  NAND2_X2 U4489 ( .A1(b[8]), .A2(a[19]), .ZN(net213477) );
  INV_X4 U4490 ( .A(net213477), .ZN(net213479) );
  INV_X32 U4491 ( .A(b[8]), .ZN(net218514) );
  NAND2_X4 U4492 ( .A1(net213479), .A2(net213478), .ZN(net213176) );
  NAND2_X2 U4493 ( .A1(net213537), .A2(net213539), .ZN(n3439) );
  XNOR2_X2 U4494 ( .A(net213538), .B(n3439), .ZN(net213787) );
  OAI21_X4 U4495 ( .B1(net212389), .B2(net219445), .A(net212413), .ZN(
        net212397) );
  XNOR2_X2 U4496 ( .A(net212122), .B(net212430), .ZN(net219412) );
  OAI21_X2 U4497 ( .B1(net212414), .B2(net212415), .A(net212416), .ZN(
        net212390) );
  INV_X4 U4498 ( .A(net212694), .ZN(net212414) );
  OAI21_X2 U4499 ( .B1(net212414), .B2(net212415), .A(net212416), .ZN(
        net219445) );
  OAI21_X4 U4500 ( .B1(net212431), .B2(net212432), .A(net220011), .ZN(
        net212122) );
  XNOR2_X2 U4501 ( .A(net212122), .B(net212394), .ZN(net212392) );
  OAI21_X2 U4502 ( .B1(net212431), .B2(net212432), .A(net220011), .ZN(
        net220298) );
  INV_X8 U4503 ( .A(net212419), .ZN(net212432) );
  XOR2_X2 U4504 ( .A(net212698), .B(net212432), .Z(net223484) );
  XNOR2_X2 U4505 ( .A(net223505), .B(net212432), .ZN(net212693) );
  INV_X1 U4506 ( .A(net220061), .ZN(net212431) );
  XNOR2_X2 U4507 ( .A(net212433), .B(n3440), .ZN(net212430) );
  XNOR2_X2 U4508 ( .A(net212430), .B(net220298), .ZN(net212389) );
  XNOR2_X2 U4509 ( .A(net212128), .B(net212393), .ZN(n3440) );
  XNOR2_X2 U4510 ( .A(net212423), .B(net212419), .ZN(net212415) );
  NAND2_X2 U4511 ( .A1(n3331), .A2(net212418), .ZN(net212416) );
  NAND2_X2 U4512 ( .A1(n3441), .A2(net213812), .ZN(net213809) );
  INV_X2 U4513 ( .A(net213810), .ZN(net213812) );
  NAND2_X2 U4514 ( .A1(a[22]), .A2(b[4]), .ZN(n3441) );
  XNOR2_X2 U4515 ( .A(net213520), .B(net213813), .ZN(net213810) );
  NAND3_X2 U4516 ( .A1(net213810), .A2(a[22]), .A3(b[4]), .ZN(net213524) );
  NAND2_X2 U4517 ( .A1(net213519), .A2(net213521), .ZN(net213813) );
  INV_X32 U4518 ( .A(b[4]), .ZN(net218530) );
  INV_X4 U4519 ( .A(net213520), .ZN(net213518) );
  OAI21_X4 U4520 ( .B1(net213517), .B2(net213518), .A(net213519), .ZN(
        net213142) );
  INV_X4 U4521 ( .A(net213521), .ZN(net213517) );
  NAND2_X4 U4522 ( .A1(n3443), .A2(net217138), .ZN(n3442) );
  OAI211_X4 U4523 ( .C1(net217127), .C2(n3442), .A(n3341), .B(net217130), .ZN(
        net217124) );
  INV_X8 U4524 ( .A(n3446), .ZN(net217138) );
  NAND3_X1 U4525 ( .A1(net217275), .A2(net217276), .A3(net217138), .ZN(
        net217274) );
  AOI21_X4 U4526 ( .B1(net217275), .B2(net217138), .A(net217278), .ZN(
        net219569) );
  NAND2_X4 U4527 ( .A1(net218081), .A2(net218082), .ZN(n3446) );
  INV_X8 U4528 ( .A(net218083), .ZN(net218081) );
  NOR2_X4 U4529 ( .A1(net217139), .A2(net217135), .ZN(n3443) );
  NAND2_X4 U4530 ( .A1(net218165), .A2(net218089), .ZN(net218082) );
  OAI21_X4 U4531 ( .B1(net217140), .B2(net218164), .A(net218082), .ZN(
        net218158) );
  NAND2_X4 U4532 ( .A1(net217136), .A2(net218159), .ZN(net218083) );
  INV_X1 U4533 ( .A(net218083), .ZN(net241365) );
  NAND2_X2 U4534 ( .A1(net218160), .A2(net218161), .ZN(net218159) );
  NAND2_X1 U4535 ( .A1(net218558), .A2(a[7]), .ZN(net218160) );
  INV_X32 U4536 ( .A(a[7]), .ZN(net218442) );
  INV_X32 U4537 ( .A(net218568), .ZN(net218558) );
  INV_X32 U4538 ( .A(b[1]), .ZN(net218568) );
  NOR2_X4 U4539 ( .A1(a[31]), .A2(net218568), .ZN(net212284) );
  INV_X32 U4540 ( .A(net218568), .ZN(net218556) );
  XNOR2_X2 U4541 ( .A(net217899), .B(net216885), .ZN(net217139) );
  OAI22_X4 U4542 ( .A1(net217139), .A2(net219569), .B1(net217276), .B2(
        net218079), .ZN(net218076) );
  INV_X4 U4543 ( .A(net217139), .ZN(net217276) );
  NAND2_X4 U4544 ( .A1(net217133), .A2(n3444), .ZN(net217135) );
  INV_X1 U4545 ( .A(net217135), .ZN(net241371) );
  NAND2_X1 U4546 ( .A1(net218558), .A2(a[9]), .ZN(n3445) );
  NAND2_X4 U4547 ( .A1(net218574), .A2(a[8]), .ZN(net218161) );
  XNOR2_X2 U4548 ( .A(net217979), .B(net218434), .ZN(net217584) );
  OAI21_X4 U4549 ( .B1(net218434), .B2(net218554), .A(net217267), .ZN(
        net216811) );
  INV_X32 U4550 ( .A(net218578), .ZN(net218574) );
  INV_X32 U4551 ( .A(b[0]), .ZN(net218578) );
  NAND2_X2 U4552 ( .A1(net218558), .A2(net218578), .ZN(net217759) );
  INV_X32 U4553 ( .A(net218578), .ZN(net218576) );
  INV_X1 U4554 ( .A(net218165), .ZN(net218224) );
  NAND3_X2 U4555 ( .A1(net218089), .A2(net218090), .A3(net218091), .ZN(
        net217141) );
  NAND2_X2 U4556 ( .A1(net218166), .A2(net218089), .ZN(net218164) );
  INV_X1 U4557 ( .A(net217136), .ZN(net217278) );
  NAND2_X2 U4558 ( .A1(a[12]), .A2(b[15]), .ZN(net213426) );
  NAND2_X4 U4559 ( .A1(net213211), .A2(net213213), .ZN(net213429) );
  OAI21_X4 U4560 ( .B1(n3447), .B2(n3448), .A(net223487), .ZN(net213212) );
  CLKBUF_X3 U4561 ( .A(net213565), .Z(net223487) );
  INV_X4 U4562 ( .A(net213567), .ZN(n3447) );
  NAND2_X4 U4563 ( .A1(net213565), .A2(net213567), .ZN(n3449) );
  XNOR2_X2 U4564 ( .A(net213566), .B(n3449), .ZN(net213745) );
  NAND2_X4 U4565 ( .A1(net213430), .A2(net213431), .ZN(net213213) );
  INV_X4 U4566 ( .A(net219990), .ZN(net213430) );
  NAND2_X2 U4567 ( .A1(a[13]), .A2(b[14]), .ZN(net213431) );
  INV_X4 U4568 ( .A(net213431), .ZN(net213433) );
  OAI22_X2 U4569 ( .A1(net216520), .A2(net218400), .B1(net216522), .B2(
        net216523), .ZN(net216334) );
  XNOR2_X2 U4570 ( .A(net216520), .B(net218400), .ZN(net216523) );
  XNOR2_X2 U4571 ( .A(net213434), .B(net213435), .ZN(net219990) );
  NAND2_X2 U4572 ( .A1(net219990), .A2(net213433), .ZN(net213211) );
  NAND2_X2 U4573 ( .A1(net213207), .A2(net213208), .ZN(net213435) );
  NAND2_X2 U4574 ( .A1(net213206), .A2(net213203), .ZN(net213434) );
  INV_X4 U4575 ( .A(net213207), .ZN(net213205) );
  NAND2_X2 U4576 ( .A1(net213750), .A2(net213208), .ZN(net213749) );
  NAND4_X2 U4577 ( .A1(a[12]), .A2(net213750), .A3(b[14]), .A4(net213208), 
        .ZN(net213565) );
  OAI21_X4 U4578 ( .B1(net213204), .B2(net213205), .A(net213206), .ZN(
        net213202) );
  NAND2_X4 U4579 ( .A1(net213202), .A2(net213203), .ZN(net212902) );
  NAND2_X4 U4580 ( .A1(net214096), .A2(net214095), .ZN(net213834) );
  OAI21_X4 U4581 ( .B1(net213833), .B2(net213311), .A(net213834), .ZN(
        net213832) );
  OAI21_X2 U4582 ( .B1(net214096), .B2(net214095), .A(net213834), .ZN(
        net214092) );
  INV_X4 U4583 ( .A(net214097), .ZN(net214096) );
  OAI21_X4 U4584 ( .B1(net214098), .B2(n3450), .A(net214100), .ZN(net214095)
         );
  INV_X8 U4585 ( .A(net214393), .ZN(net214098) );
  XNOR2_X2 U4586 ( .A(net214098), .B(n3451), .ZN(net214385) );
  OAI21_X4 U4587 ( .B1(net214394), .B2(net213634), .A(net214395), .ZN(
        net214393) );
  XNOR2_X2 U4588 ( .A(net213833), .B(net213311), .ZN(net214097) );
  INV_X4 U4589 ( .A(n3450), .ZN(n3451) );
  NAND2_X2 U4590 ( .A1(net214100), .A2(net214389), .ZN(n3450) );
  XNOR2_X2 U4591 ( .A(net214394), .B(net213634), .ZN(net214665) );
  NAND2_X4 U4592 ( .A1(net216068), .A2(net216067), .ZN(net215856) );
  OAI21_X4 U4593 ( .B1(net215855), .B2(net215245), .A(net215856), .ZN(
        net215854) );
  OAI21_X2 U4594 ( .B1(net216068), .B2(net219557), .A(net215856), .ZN(
        net216064) );
  INV_X4 U4595 ( .A(net216069), .ZN(net216068) );
  OAI21_X4 U4596 ( .B1(net216070), .B2(n3452), .A(net216072), .ZN(net216067)
         );
  XNOR2_X2 U4597 ( .A(net215855), .B(net215245), .ZN(net216069) );
  XNOR2_X2 U4598 ( .A(net216252), .B(n3452), .ZN(net216052) );
  NAND2_X2 U4599 ( .A1(net216253), .A2(net216072), .ZN(n3452) );
  NAND2_X2 U4600 ( .A1(n3454), .A2(net216965), .ZN(net216962) );
  NAND2_X2 U4601 ( .A1(net218558), .A2(a[11]), .ZN(n3454) );
  OAI22_X2 U4602 ( .A1(net216998), .A2(net218414), .B1(net217000), .B2(
        net217001), .ZN(net216716) );
  XNOR2_X2 U4603 ( .A(net216998), .B(net218414), .ZN(net217001) );
  NAND2_X2 U4604 ( .A1(n3453), .A2(a[11]), .ZN(net216800) );
  INV_X4 U4605 ( .A(net216328), .ZN(n3453) );
  NAND2_X4 U4606 ( .A1(net213447), .A2(net213446), .ZN(net213206) );
  INV_X4 U4607 ( .A(net213445), .ZN(net213447) );
  XNOR2_X2 U4608 ( .A(net213448), .B(net213449), .ZN(net213445) );
  NAND2_X2 U4609 ( .A1(net213444), .A2(net224038), .ZN(net213203) );
  XNOR2_X2 U4610 ( .A(net213448), .B(net213449), .ZN(net224038) );
  INV_X4 U4611 ( .A(net213446), .ZN(net213444) );
  NAND2_X2 U4612 ( .A1(a[11]), .A2(b[16]), .ZN(net213421) );
  INV_X4 U4613 ( .A(net213217), .ZN(net213215) );
  NAND2_X2 U4614 ( .A1(a[9]), .A2(b[19]), .ZN(net213045) );
  NAND2_X2 U4615 ( .A1(a[10]), .A2(b[18]), .ZN(net213050) );
  NAND2_X4 U4616 ( .A1(net212920), .A2(net212921), .ZN(net213054) );
  INV_X2 U4617 ( .A(net212921), .ZN(net212918) );
  XNOR2_X2 U4618 ( .A(net213414), .B(net213413), .ZN(net213411) );
  NOR2_X4 U4619 ( .A1(net223606), .A2(net223578), .ZN(net223577) );
  INV_X2 U4620 ( .A(net223577), .ZN(net211934) );
  NOR3_X2 U4621 ( .A1(net211942), .A2(net223577), .A3(net211944), .ZN(zero) );
  INV_X32 U4622 ( .A(net218658), .ZN(net218660) );
  NAND3_X4 U4623 ( .A1(op[2]), .A2(op[0]), .A3(n3455), .ZN(net212100) );
  INV_X4 U4624 ( .A(n3458), .ZN(n3455) );
  NAND3_X4 U4625 ( .A1(n3455), .A2(net217946), .A3(net217346), .ZN(net211949)
         );
  NAND3_X4 U4626 ( .A1(op[0]), .A2(n3455), .A3(net217946), .ZN(net211950) );
  NAND2_X2 U4627 ( .A1(n3456), .A2(n3457), .ZN(n3458) );
  INV_X4 U4628 ( .A(op[1]), .ZN(n3457) );
  INV_X4 U4629 ( .A(op[3]), .ZN(n3456) );
  NAND2_X2 U4630 ( .A1(op[1]), .A2(n3456), .ZN(net217948) );
  XNOR2_X2 U4631 ( .A(net212104), .B(net223607), .ZN(net223606) );
  XNOR2_X2 U4632 ( .A(net212110), .B(net212111), .ZN(net223607) );
  INV_X4 U4633 ( .A(b[31]), .ZN(net212023) );
  NAND2_X2 U4634 ( .A1(b[31]), .A2(net217557), .ZN(net217362) );
  NAND2_X4 U4635 ( .A1(net218658), .A2(net218496), .ZN(net212094) );
  INV_X4 U4636 ( .A(a[0]), .ZN(net218496) );
  NAND2_X2 U4637 ( .A1(op[3]), .A2(net217348), .ZN(net217340) );
  NAND2_X2 U4638 ( .A1(op[3]), .A2(op[2]), .ZN(net217966) );
  INV_X4 U4639 ( .A(op[3]), .ZN(net218370) );
  NAND2_X4 U4640 ( .A1(net223109), .A2(net212105), .ZN(net212104) );
  XNOR2_X2 U4641 ( .A(net212103), .B(net212104), .ZN(net212099) );
  NAND2_X4 U4642 ( .A1(net212934), .A2(net212936), .ZN(net213038) );
  NAND2_X2 U4643 ( .A1(net213042), .A2(net213041), .ZN(net212934) );
  INV_X4 U4644 ( .A(net213040), .ZN(net213042) );
  NAND2_X4 U4645 ( .A1(net213039), .A2(net213040), .ZN(net212936) );
  INV_X2 U4646 ( .A(net212936), .ZN(net212932) );
  INV_X4 U4647 ( .A(net213041), .ZN(net213039) );
  INV_X4 U4648 ( .A(net215184), .ZN(net215181) );
  NAND2_X4 U4649 ( .A1(n3459), .A2(net215640), .ZN(net215185) );
  OAI21_X2 U4650 ( .B1(net215640), .B2(net220060), .A(net215185), .ZN(
        net215636) );
  INV_X4 U4651 ( .A(net215641), .ZN(net215640) );
  OAI21_X4 U4652 ( .B1(net215642), .B2(net215643), .A(net215644), .ZN(n3459)
         );
  INV_X8 U4653 ( .A(net215854), .ZN(net215642) );
  OAI21_X1 U4654 ( .B1(net215642), .B2(net215643), .A(net215644), .ZN(
        net220060) );
  XNOR2_X2 U4655 ( .A(net215642), .B(net215849), .ZN(net215846) );
  NAND2_X2 U4656 ( .A1(net215422), .A2(net215423), .ZN(net215186) );
  INV_X4 U4657 ( .A(net215424), .ZN(net215423) );
  INV_X4 U4658 ( .A(net215001), .ZN(net215422) );
  INV_X4 U4659 ( .A(net215643), .ZN(net215849) );
  NAND2_X2 U4660 ( .A1(net215850), .A2(net215644), .ZN(net215643) );
  XNOR2_X2 U4661 ( .A(net215424), .B(net215001), .ZN(net215641) );
  INV_X4 U4662 ( .A(b[30]), .ZN(n3460) );
  NAND2_X2 U4663 ( .A1(net218658), .A2(n3460), .ZN(net212093) );
  INV_X4 U4664 ( .A(net223126), .ZN(net223109) );
  AND2_X2 U4665 ( .A1(net223109), .A2(net212092), .ZN(net223617) );
  NOR2_X1 U4666 ( .A1(net218655), .A2(net223109), .ZN(net211946) );
  XNOR2_X2 U4667 ( .A(net223104), .B(net223100), .ZN(net223126) );
  XNOR2_X2 U4668 ( .A(net223498), .B(net223124), .ZN(net223481) );
  XNOR2_X2 U4669 ( .A(net212405), .B(net212402), .ZN(net223125) );
  XNOR2_X2 U4670 ( .A(net212405), .B(net212402), .ZN(net223498) );
  NAND3_X4 U4671 ( .A1(b[29]), .A2(a[0]), .A3(net223098), .ZN(net223100) );
  OAI21_X4 U4672 ( .B1(net223100), .B2(net223481), .A(net223105), .ZN(
        net212110) );
  INV_X8 U4673 ( .A(net212672), .ZN(net223098) );
  OAI21_X4 U4674 ( .B1(net218655), .B2(net223098), .A(net212681), .ZN(
        net212679) );
  NAND2_X4 U4675 ( .A1(net212403), .A2(n3429), .ZN(net223009) );
  XNOR2_X2 U4676 ( .A(net212399), .B(net223009), .ZN(net212401) );
  NAND2_X2 U4677 ( .A1(n3461), .A2(net212411), .ZN(net212403) );
  INV_X4 U4678 ( .A(net212412), .ZN(n3461) );
  NAND2_X4 U4679 ( .A1(net223089), .A2(net223090), .ZN(net212405) );
  INV_X2 U4680 ( .A(net212405), .ZN(net212399) );
  NAND2_X4 U4681 ( .A1(net213198), .A2(net212794), .ZN(net213449) );
  NAND2_X2 U4682 ( .A1(net213453), .A2(net213452), .ZN(net213198) );
  NAND2_X2 U4683 ( .A1(net213197), .A2(net213198), .ZN(net212795) );
  INV_X2 U4684 ( .A(net213451), .ZN(net213453) );
  NAND3_X1 U4685 ( .A1(net212794), .A2(net212636), .A3(net212795), .ZN(
        net212792) );
  INV_X4 U4686 ( .A(net213452), .ZN(net213450) );
  NAND2_X2 U4687 ( .A1(net213182), .A2(net213184), .ZN(net213466) );
  XNOR2_X2 U4688 ( .A(net213183), .B(net213466), .ZN(net213463) );
  NAND2_X2 U4689 ( .A1(net213470), .A2(net213469), .ZN(net213182) );
  OAI21_X4 U4690 ( .B1(net213180), .B2(net213181), .A(net213182), .ZN(
        net212888) );
  INV_X4 U4691 ( .A(net213468), .ZN(net213470) );
  NAND2_X2 U4692 ( .A1(net213467), .A2(net213468), .ZN(net213184) );
  INV_X4 U4693 ( .A(net213184), .ZN(net213180) );
  INV_X4 U4694 ( .A(net213469), .ZN(net213467) );
  NAND3_X2 U4695 ( .A1(a[23]), .A2(net213816), .A3(net218534), .ZN(net213519)
         );
  INV_X32 U4696 ( .A(net218544), .ZN(net218534) );
  INV_X32 U4697 ( .A(b[3]), .ZN(net218544) );
  INV_X4 U4698 ( .A(net220036), .ZN(net213816) );
  NAND2_X2 U4699 ( .A1(net213814), .A2(net220036), .ZN(net213521) );
  NAND2_X2 U4700 ( .A1(a[23]), .A2(net218538), .ZN(net213814) );
  INV_X32 U4701 ( .A(net218542), .ZN(net218538) );
  INV_X32 U4702 ( .A(b[3]), .ZN(net218542) );
  INV_X32 U4703 ( .A(net218542), .ZN(net218536) );
  NAND2_X2 U4704 ( .A1(net213166), .A2(net213168), .ZN(net213490) );
  XNOR2_X2 U4705 ( .A(net213167), .B(net213490), .ZN(net213488) );
  NAND2_X2 U4706 ( .A1(net213494), .A2(net213493), .ZN(net213166) );
  OAI21_X4 U4707 ( .B1(net213164), .B2(net213165), .A(net213166), .ZN(
        net212842) );
  INV_X4 U4708 ( .A(net213491), .ZN(net213494) );
  INV_X4 U4709 ( .A(net213168), .ZN(net213164) );
  INV_X4 U4710 ( .A(net213493), .ZN(net213492) );
  NAND2_X2 U4711 ( .A1(net213114), .A2(net213116), .ZN(net213485) );
  XNOR2_X2 U4712 ( .A(net213115), .B(net213485), .ZN(net213483) );
  NAND2_X2 U4713 ( .A1(net213489), .A2(net213488), .ZN(net213114) );
  OAI21_X4 U4714 ( .B1(net213112), .B2(net213113), .A(net213114), .ZN(
        net213111) );
  INV_X4 U4715 ( .A(net213486), .ZN(net213489) );
  NAND2_X2 U4716 ( .A1(net213486), .A2(net213487), .ZN(net213116) );
  INV_X4 U4717 ( .A(net213116), .ZN(net213112) );
  INV_X4 U4718 ( .A(net213488), .ZN(net213487) );
  NAND2_X2 U4719 ( .A1(net213484), .A2(net213483), .ZN(net213171) );
  INV_X4 U4720 ( .A(net213481), .ZN(net213484) );
  NAND2_X2 U4721 ( .A1(net213481), .A2(net213482), .ZN(net213173) );
  INV_X4 U4722 ( .A(net213483), .ZN(net213482) );
  NAND2_X2 U4723 ( .A1(net213189), .A2(net213186), .ZN(net213461) );
  XNOR2_X2 U4724 ( .A(net213460), .B(net213461), .ZN(net213457) );
  NAND2_X4 U4725 ( .A1(net213465), .A2(net213464), .ZN(net213189) );
  OAI21_X4 U4726 ( .B1(net213187), .B2(net213188), .A(net213189), .ZN(
        net213185) );
  INV_X4 U4727 ( .A(net213463), .ZN(net213465) );
  NAND2_X2 U4728 ( .A1(net213462), .A2(net213463), .ZN(net213186) );
  NAND2_X4 U4729 ( .A1(net213185), .A2(net213186), .ZN(net212893) );
  INV_X4 U4730 ( .A(net213464), .ZN(net213462) );
  NAND2_X2 U4731 ( .A1(n3463), .A2(net215853), .ZN(net215850) );
  NAND2_X2 U4732 ( .A1(net218556), .A2(a[17]), .ZN(n3463) );
  INV_X32 U4733 ( .A(a[17]), .ZN(net218378) );
  NAND2_X2 U4734 ( .A1(n3462), .A2(a[17]), .ZN(net215644) );
  INV_X4 U4735 ( .A(net215023), .ZN(n3462) );
  NAND2_X2 U4736 ( .A1(net218574), .A2(a[17]), .ZN(net215245) );
  NAND4_X1 U4737 ( .A1(net217027), .A2(net217028), .A3(net217029), .A4(
        net217030), .ZN(net214477) );
  NAND4_X1 U4738 ( .A1(net217859), .A2(net217028), .A3(net217860), .A4(
        net217621), .ZN(net217858) );
  NAND2_X1 U4739 ( .A1(net217970), .A2(net218566), .ZN(net217816) );
  NAND2_X4 U4740 ( .A1(net215177), .A2(net215178), .ZN(net214930) );
  OAI21_X4 U4741 ( .B1(net214929), .B2(net214224), .A(net214930), .ZN(
        net214928) );
  OAI21_X4 U4742 ( .B1(net215181), .B2(n3464), .A(net215183), .ZN(net215178)
         );
  XNOR2_X2 U4743 ( .A(net214929), .B(net214224), .ZN(net215180) );
  INV_X4 U4744 ( .A(net215180), .ZN(net215177) );
  XNOR2_X2 U4745 ( .A(net215417), .B(n3464), .ZN(net215414) );
  NAND2_X2 U4746 ( .A1(net215418), .A2(net215183), .ZN(n3464) );
  NAND2_X4 U4747 ( .A1(net214662), .A2(net214663), .ZN(net214395) );
  OAI21_X4 U4748 ( .B1(net214666), .B2(n3465), .A(net214668), .ZN(net214663)
         );
  INV_X8 U4749 ( .A(net214928), .ZN(net214666) );
  XNOR2_X2 U4750 ( .A(net214666), .B(n3466), .ZN(net214922) );
  INV_X4 U4751 ( .A(net214665), .ZN(net214662) );
  INV_X4 U4752 ( .A(n3465), .ZN(n3466) );
  NAND2_X2 U4753 ( .A1(net214668), .A2(net214924), .ZN(n3465) );
  NAND2_X2 U4754 ( .A1(n3467), .A2(net211939), .ZN(net211944) );
  NOR3_X2 U4755 ( .A1(net223617), .A2(n7897), .A3(n3306), .ZN(n3467) );
  NAND2_X2 U4756 ( .A1(n3469), .A2(n3470), .ZN(n3468) );
  INV_X4 U4757 ( .A(result[17]), .ZN(n3470) );
  NOR2_X4 U4758 ( .A1(result[16]), .A2(n3351), .ZN(n3469) );
  NAND2_X4 U4759 ( .A1(net213016), .A2(net213015), .ZN(net212946) );
  NAND2_X4 U4760 ( .A1(net212944), .A2(net212946), .ZN(net213012) );
  INV_X4 U4761 ( .A(net212946), .ZN(net212945) );
  INV_X4 U4762 ( .A(net213013), .ZN(net213016) );
  INV_X4 U4763 ( .A(net213014), .ZN(net213015) );
  NAND2_X2 U4764 ( .A1(net213014), .A2(net213013), .ZN(net212944) );
  NAND3_X2 U4765 ( .A1(net213021), .A2(net213384), .A3(net220146), .ZN(
        net213020) );
  INV_X4 U4766 ( .A(net220145), .ZN(net220146) );
  NAND2_X4 U4767 ( .A1(net213021), .A2(net220146), .ZN(net212735) );
  INV_X2 U4768 ( .A(net213022), .ZN(net220145) );
  NAND2_X2 U4769 ( .A1(a[5]), .A2(b[23]), .ZN(net213014) );
  NAND2_X4 U4770 ( .A1(net213608), .A2(net213022), .ZN(net213692) );
  NAND2_X4 U4771 ( .A1(net213823), .A2(net213516), .ZN(net213515) );
  OAI21_X4 U4772 ( .B1(net213514), .B2(net213515), .A(net223812), .ZN(
        net213152) );
  XNOR2_X2 U4773 ( .A(net213515), .B(net213514), .ZN(net220036) );
  NAND2_X2 U4774 ( .A1(n3471), .A2(net213826), .ZN(net213823) );
  INV_X4 U4775 ( .A(net213824), .ZN(net213826) );
  NAND2_X2 U4776 ( .A1(a[24]), .A2(net218550), .ZN(n3471) );
  INV_X32 U4777 ( .A(net218552), .ZN(net218550) );
  INV_X32 U4778 ( .A(b[2]), .ZN(net218552) );
  INV_X32 U4779 ( .A(net218552), .ZN(net218546) );
  INV_X32 U4780 ( .A(net218552), .ZN(net218548) );
  NAND3_X2 U4781 ( .A1(a[24]), .A2(net213824), .A3(net218548), .ZN(net213516)
         );
  CLKBUF_X3 U4782 ( .A(net213516), .Z(net223812) );
  XNOR2_X2 U4783 ( .A(net213511), .B(n3472), .ZN(net213824) );
  INV_X4 U4784 ( .A(net213512), .ZN(n3472) );
  INV_X4 U4785 ( .A(net213832), .ZN(net213511) );
  OAI21_X4 U4786 ( .B1(net213511), .B2(net213512), .A(net213513), .ZN(
        net213508) );
  INV_X32 U4787 ( .A(b[2]), .ZN(net218554) );
  NOR2_X4 U4788 ( .A1(net217131), .A2(n3473), .ZN(net217130) );
  INV_X4 U4789 ( .A(n3474), .ZN(n3473) );
  NOR2_X2 U4790 ( .A1(net217278), .A2(n3473), .ZN(net217273) );
  NAND2_X2 U4791 ( .A1(net217183), .A2(net217280), .ZN(n3474) );
  INV_X4 U4792 ( .A(net217899), .ZN(net217280) );
  NAND2_X2 U4793 ( .A1(net217280), .A2(net218578), .ZN(net217182) );
  INV_X4 U4794 ( .A(net216885), .ZN(net217183) );
  NAND2_X2 U4795 ( .A1(net217183), .A2(net218566), .ZN(net217179) );
  INV_X4 U4796 ( .A(net217133), .ZN(net217131) );
  INV_X8 U4797 ( .A(net217142), .ZN(net217140) );
  NAND2_X4 U4798 ( .A1(n3300), .A2(a[7]), .ZN(net217136) );
  NAND2_X4 U4799 ( .A1(net212722), .A2(net212721), .ZN(net212647) );
  INV_X4 U4800 ( .A(net212720), .ZN(net212722) );
  NAND2_X2 U4801 ( .A1(b[24]), .A2(a[5]), .ZN(net212721) );
  INV_X4 U4802 ( .A(net212721), .ZN(net212719) );
  XNOR2_X2 U4803 ( .A(net212723), .B(net212724), .ZN(net212720) );
  NAND2_X2 U4804 ( .A1(net212719), .A2(net212720), .ZN(net212648) );
  NAND2_X2 U4805 ( .A1(net212454), .A2(n3477), .ZN(net212724) );
  NAND2_X2 U4806 ( .A1(net241088), .A2(net241082), .ZN(n3477) );
  INV_X4 U4807 ( .A(n3475), .ZN(net212723) );
  AOI21_X4 U4808 ( .B1(n3476), .B2(net212944), .A(net212945), .ZN(n3475) );
  OAI21_X1 U4809 ( .B1(net212452), .B2(n3475), .A(net212454), .ZN(net212451)
         );
  INV_X4 U4810 ( .A(net241082), .ZN(net241076) );
  NAND2_X4 U4811 ( .A1(net213250), .A2(net212948), .ZN(net213381) );
  NAND2_X2 U4812 ( .A1(net212397), .A2(net212398), .ZN(net223090) );
  INV_X4 U4813 ( .A(net212397), .ZN(net223121) );
  NAND2_X2 U4814 ( .A1(b[28]), .A2(a[2]), .ZN(net212398) );
  INV_X4 U4815 ( .A(net212398), .ZN(net223119) );
  NAND2_X1 U4816 ( .A1(net217654), .A2(net218476), .ZN(net218353) );
  XNOR2_X1 U4817 ( .A(net217995), .B(net218476), .ZN(net217933) );
  NAND2_X1 U4818 ( .A1(net218548), .A2(net218476), .ZN(net217431) );
  NAND2_X4 U4819 ( .A1(net223121), .A2(net223119), .ZN(net223089) );
  NAND2_X1 U4820 ( .A1(net223119), .A2(net223121), .ZN(net223586) );
  NAND2_X2 U4821 ( .A1(a[24]), .A2(net218556), .ZN(net213833) );
  NAND2_X2 U4822 ( .A1(a[25]), .A2(net218576), .ZN(net213311) );
  INV_X4 U4823 ( .A(net216965), .ZN(net217818) );
  NAND4_X2 U4824 ( .A1(net216327), .A2(net216328), .A3(net216329), .A4(
        net216330), .ZN(net213359) );
  INV_X4 U4825 ( .A(net215853), .ZN(net217807) );
  OAI21_X4 U4826 ( .B1(net216444), .B2(n3478), .A(net216446), .ZN(net216441)
         );
  XNOR2_X2 U4827 ( .A(net216623), .B(n3478), .ZN(net216620) );
  NAND2_X2 U4828 ( .A1(net216624), .A2(net216446), .ZN(n3478) );
  NAND2_X2 U4829 ( .A1(a[7]), .A2(b[21]), .ZN(net213036) );
  OAI21_X4 U4830 ( .B1(net213241), .B2(net213240), .A(n3199), .ZN(net212935)
         );
  INV_X2 U4831 ( .A(net213248), .ZN(net213240) );
  AOI21_X2 U4832 ( .B1(net213243), .B2(net213244), .A(net213245), .ZN(
        net213241) );
  INV_X1 U4833 ( .A(net213245), .ZN(net220046) );
  NOR2_X4 U4834 ( .A1(net213247), .A2(net213245), .ZN(net213700) );
  NOR3_X2 U4835 ( .A1(n3302), .A2(net213603), .A3(net213245), .ZN(net213704)
         );
  NAND2_X2 U4836 ( .A1(net213711), .A2(n3479), .ZN(net213596) );
  INV_X4 U4837 ( .A(net213712), .ZN(n3479) );
  NOR2_X2 U4838 ( .A1(n3302), .A2(net213246), .ZN(net213243) );
  AOI21_X4 U4839 ( .B1(net213702), .B2(net213703), .A(net213246), .ZN(
        net213701) );
  NAND2_X4 U4840 ( .A1(net213242), .A2(net213248), .ZN(net213398) );
  OAI21_X4 U4841 ( .B1(n3480), .B2(n3207), .A(net213201), .ZN(net213448) );
  OAI21_X2 U4842 ( .B1(n3480), .B2(n3207), .A(net213201), .ZN(net213197) );
  OAI21_X2 U4843 ( .B1(net213560), .B2(net213870), .A(net213562), .ZN(n3482)
         );
  OAI21_X4 U4844 ( .B1(net214326), .B2(net213870), .A(net214325), .ZN(
        net214152) );
  INV_X4 U4845 ( .A(net213442), .ZN(n3480) );
  NAND2_X2 U4846 ( .A1(net213201), .A2(net213442), .ZN(net213438) );
  NAND2_X4 U4847 ( .A1(n3481), .A2(net213441), .ZN(net213439) );
  NAND2_X2 U4848 ( .A1(net213441), .A2(net213562), .ZN(net214019) );
  NOR2_X4 U4849 ( .A1(net213870), .A2(net213560), .ZN(net214020) );
  NAND3_X2 U4850 ( .A1(net214323), .A2(net214025), .A3(net214324), .ZN(
        net214147) );
  NAND2_X4 U4851 ( .A1(net213249), .A2(net213250), .ZN(net212947) );
  NAND2_X4 U4852 ( .A1(net213251), .A2(net219874), .ZN(net213249) );
  NAND2_X4 U4853 ( .A1(net213386), .A2(n3483), .ZN(net212948) );
  XNOR2_X2 U4854 ( .A(net212735), .B(n3244), .ZN(net213386) );
  INV_X4 U4855 ( .A(net213383), .ZN(n3483) );
  NAND2_X2 U4856 ( .A1(net219874), .A2(net213251), .ZN(net213380) );
  XNOR2_X2 U4857 ( .A(n3244), .B(net212732), .ZN(net213382) );
  NAND2_X4 U4858 ( .A1(net213382), .A2(net213383), .ZN(net213250) );
  NAND2_X2 U4859 ( .A1(a[22]), .A2(b[5]), .ZN(net213491) );
  XNOR2_X2 U4860 ( .A(net213131), .B(net213495), .ZN(net213493) );
  INV_X4 U4861 ( .A(net213131), .ZN(net213129) );
  OAI21_X2 U4862 ( .B1(n3484), .B2(net213129), .A(net213130), .ZN(net213127)
         );
  NAND2_X2 U4863 ( .A1(a[21]), .A2(b[6]), .ZN(net213486) );
  NAND2_X2 U4864 ( .A1(a[6]), .A2(n3485), .ZN(net217524) );
  NOR2_X4 U4865 ( .A1(a[6]), .A2(n3485), .ZN(net217438) );
  INV_X4 U4866 ( .A(net213167), .ZN(net213165) );
  NAND2_X2 U4867 ( .A1(b[7]), .A2(a[20]), .ZN(net213481) );
  INV_X4 U4868 ( .A(net213115), .ZN(net213113) );
  NAND2_X2 U4869 ( .A1(net218556), .A2(a[20]), .ZN(net214929) );
  NAND2_X2 U4870 ( .A1(a[21]), .A2(net218576), .ZN(net214224) );
  NAND2_X2 U4871 ( .A1(a[22]), .A2(net218558), .ZN(net214394) );
  NAND2_X2 U4872 ( .A1(a[23]), .A2(net218576), .ZN(net213634) );
  NAND2_X2 U4873 ( .A1(net213190), .A2(net213191), .ZN(net213460) );
  NAND2_X2 U4874 ( .A1(a[16]), .A2(b[11]), .ZN(net213458) );
  NAND2_X2 U4875 ( .A1(a[11]), .A2(n3486), .ZN(net217512) );
  NOR2_X4 U4876 ( .A1(a[11]), .A2(n3486), .ZN(net217414) );
  INV_X4 U4877 ( .A(net213190), .ZN(net213188) );
  INV_X2 U4878 ( .A(net213191), .ZN(net213187) );
  NAND2_X2 U4879 ( .A1(net213546), .A2(net213191), .ZN(net213773) );
  NAND2_X2 U4880 ( .A1(b[25]), .A2(a[4]), .ZN(net212441) );
  NAND3_X2 U4881 ( .A1(b[4]), .A2(net217445), .A3(net219068), .ZN(net217442)
         );
  NAND2_X2 U4882 ( .A1(net213418), .A2(net213417), .ZN(net213227) );
  INV_X4 U4883 ( .A(net213416), .ZN(net213418) );
  NAND2_X2 U4884 ( .A1(a[10]), .A2(b[17]), .ZN(net213416) );
  NAND2_X4 U4885 ( .A1(net213415), .A2(net213416), .ZN(net213225) );
  INV_X4 U4886 ( .A(net213222), .ZN(net213220) );
  OAI21_X2 U4887 ( .B1(net213522), .B2(net213523), .A(net213524), .ZN(
        net213131) );
  INV_X4 U4888 ( .A(net213523), .ZN(net213804) );
  NAND2_X2 U4889 ( .A1(a[15]), .A2(b[12]), .ZN(net213452) );
  OAI22_X2 U4890 ( .A1(net216126), .A2(n3487), .B1(net216128), .B2(net216129), 
        .ZN(net215913) );
  XNOR2_X2 U4891 ( .A(net216126), .B(n3487), .ZN(net216129) );
  NAND2_X2 U4892 ( .A1(net213195), .A2(net213196), .ZN(net213454) );
  INV_X2 U4893 ( .A(net213195), .ZN(net213193) );
  NAND2_X2 U4894 ( .A1(net213551), .A2(net213196), .ZN(net213767) );
  NAND2_X2 U4895 ( .A1(n3489), .A2(net216256), .ZN(net216253) );
  NAND2_X2 U4896 ( .A1(net218558), .A2(a[15]), .ZN(n3489) );
  NAND2_X2 U4897 ( .A1(n3488), .A2(a[15]), .ZN(net216072) );
  INV_X4 U4898 ( .A(net215492), .ZN(n3488) );
  INV_X4 U4899 ( .A(net216256), .ZN(net217806) );
  NAND4_X2 U4900 ( .A1(net216711), .A2(net215492), .A3(net215920), .A4(
        net216327), .ZN(net216704) );
  NAND4_X2 U4901 ( .A1(net215491), .A2(net215492), .A3(net215493), .A4(
        net215494), .ZN(net212010) );
  NAND2_X2 U4902 ( .A1(a[18]), .A2(b[9]), .ZN(net213468) );
  NAND2_X2 U4903 ( .A1(b[29]), .A2(net218480), .ZN(net212402) );
  NOR2_X2 U4904 ( .A1(net212401), .A2(net212402), .ZN(net223123) );
  NAND2_X2 U4905 ( .A1(b[26]), .A2(net218480), .ZN(net213367) );
  NAND2_X2 U4906 ( .A1(b[28]), .A2(net218480), .ZN(net212688) );
  NAND2_X2 U4907 ( .A1(net212411), .A2(net212404), .ZN(net212683) );
  XNOR2_X2 U4908 ( .A(net212683), .B(net212412), .ZN(net212672) );
  NAND2_X2 U4909 ( .A1(n3491), .A2(net216627), .ZN(net216624) );
  NAND2_X2 U4910 ( .A1(a[13]), .A2(net218558), .ZN(n3491) );
  NAND2_X2 U4911 ( .A1(a[13]), .A2(n3490), .ZN(net216446) );
  INV_X4 U4912 ( .A(net215919), .ZN(n3490) );
  NAND2_X2 U4913 ( .A1(n3492), .A2(net214391), .ZN(net214389) );
  NAND2_X2 U4914 ( .A1(a[23]), .A2(net218558), .ZN(n3492) );
  NAND2_X2 U4915 ( .A1(n3493), .A2(a[23]), .ZN(net214100) );
  INV_X4 U4916 ( .A(net213331), .ZN(n3493) );
  INV_X4 U4917 ( .A(net214391), .ZN(net217783) );
  NAND4_X2 U4918 ( .A1(net214486), .A2(net213331), .A3(net213926), .A4(
        net215024), .ZN(net217838) );
  NAND4_X2 U4919 ( .A1(net213330), .A2(net213331), .A3(net213332), .A4(
        net213333), .ZN(net212007) );
  NAND2_X2 U4920 ( .A1(b[13]), .A2(a[14]), .ZN(net213446) );
  NOR2_X4 U4921 ( .A1(a[13]), .A2(net218502), .ZN(net217408) );
  NAND2_X2 U4922 ( .A1(a[13]), .A2(net218502), .ZN(net217506) );
  NAND2_X2 U4923 ( .A1(a[17]), .A2(b[10]), .ZN(net213464) );
  INV_X4 U4924 ( .A(net213183), .ZN(net213181) );
  NOR2_X4 U4925 ( .A1(net213706), .A2(net213603), .ZN(net213705) );
  NAND2_X4 U4926 ( .A1(net213602), .A2(net213603), .ZN(net213607) );
  XNOR2_X2 U4927 ( .A(net213700), .B(net213701), .ZN(net213602) );
  INV_X2 U4928 ( .A(net213244), .ZN(net213706) );
  NAND3_X2 U4929 ( .A1(net220017), .A2(net213244), .A3(n3194), .ZN(net213595)
         );
  INV_X2 U4930 ( .A(net213711), .ZN(net213713) );
  NAND2_X4 U4931 ( .A1(net213713), .A2(net213712), .ZN(net213597) );
  NAND2_X4 U4932 ( .A1(net213703), .A2(net213598), .ZN(net213969) );
  XNOR2_X2 U4933 ( .A(net212419), .B(net212420), .ZN(net212418) );
  XNOR2_X2 U4934 ( .A(net212420), .B(n3331), .ZN(net223505) );
  XNOR2_X2 U4935 ( .A(net212420), .B(n3331), .ZN(net212698) );
  NAND2_X4 U4936 ( .A1(net219338), .A2(n3363), .ZN(net212429) );
  NAND2_X2 U4937 ( .A1(a[8]), .A2(b[20]), .ZN(net213040) );
  INV_X4 U4938 ( .A(net212930), .ZN(net212928) );
  NAND2_X2 U4939 ( .A1(n3494), .A2(net213229), .ZN(net213413) );
  NAND2_X2 U4940 ( .A1(net213580), .A2(net213581), .ZN(n3494) );
  OAI21_X2 U4941 ( .B1(n3495), .B2(net213583), .A(n3502), .ZN(net213580) );
  INV_X4 U4942 ( .A(n3498), .ZN(n3502) );
  INV_X4 U4943 ( .A(n3496), .ZN(n3498) );
  NOR2_X4 U4944 ( .A1(n3501), .A2(n3498), .ZN(net213725) );
  NOR2_X4 U4945 ( .A1(n3498), .A2(n3495), .ZN(n3499) );
  NAND2_X2 U4946 ( .A1(n3500), .A2(n3503), .ZN(n3496) );
  INV_X4 U4947 ( .A(net213994), .ZN(n3500) );
  INV_X2 U4948 ( .A(net213726), .ZN(net213583) );
  XNOR2_X2 U4949 ( .A(n3499), .B(net213583), .ZN(net213984) );
  INV_X8 U4950 ( .A(n3497), .ZN(n3495) );
  NAND2_X4 U4951 ( .A1(net213229), .A2(net213581), .ZN(net213729) );
  XNOR2_X2 U4952 ( .A(net213997), .B(net213576), .ZN(net213995) );
  AOI21_X4 U4953 ( .B1(net213576), .B2(n3192), .A(net213578), .ZN(net213574)
         );
  NAND2_X4 U4954 ( .A1(net213993), .A2(net213994), .ZN(n3497) );
  AND2_X2 U4955 ( .A1(net213726), .A2(n3497), .ZN(n3501) );
  XNOR2_X2 U4956 ( .A(net212110), .B(net212111), .ZN(net212103) );
  INV_X4 U4957 ( .A(net223123), .ZN(net223105) );
  NAND2_X2 U4958 ( .A1(n3505), .A2(net215421), .ZN(net215418) );
  NAND2_X2 U4959 ( .A1(a[19]), .A2(net218558), .ZN(n3505) );
  NAND2_X2 U4960 ( .A1(a[19]), .A2(n3504), .ZN(net215183) );
  NOR2_X4 U4961 ( .A1(net215421), .A2(n3301), .ZN(n3504) );
  INV_X4 U4962 ( .A(net215421), .ZN(net217781) );
  INV_X4 U4963 ( .A(n3504), .ZN(net214487) );
  NAND2_X2 U4964 ( .A1(n3506), .A2(net214926), .ZN(net214924) );
  NAND2_X2 U4965 ( .A1(a[21]), .A2(net218556), .ZN(n3506) );
  NAND2_X2 U4966 ( .A1(n3507), .A2(a[21]), .ZN(net214668) );
  INV_X4 U4967 ( .A(net213925), .ZN(n3507) );
  INV_X4 U4968 ( .A(net214926), .ZN(net217780) );
  NAND4_X2 U4969 ( .A1(net215022), .A2(net213925), .A3(net215493), .A4(
        net214489), .ZN(net217779) );
  NAND4_X2 U4970 ( .A1(net213924), .A2(net213925), .A3(net213926), .A4(
        net213927), .ZN(net212971) );
  AOI21_X4 U4971 ( .B1(n3510), .B2(net213553), .A(n3511), .ZN(n3509) );
  NAND2_X1 U4972 ( .A1(net213556), .A2(net213557), .ZN(n3510) );
  AOI21_X2 U4973 ( .B1(net213763), .B2(net213555), .A(n3508), .ZN(net213762)
         );
  NAND2_X2 U4974 ( .A1(n3512), .A2(net213769), .ZN(net213196) );
  INV_X4 U4975 ( .A(net213770), .ZN(n3512) );
  NAND2_X4 U4976 ( .A1(net213555), .A2(net213764), .ZN(net214033) );
  INV_X4 U4977 ( .A(net213556), .ZN(net213766) );
  INV_X2 U4978 ( .A(net213769), .ZN(n3513) );
  OAI21_X4 U4979 ( .B1(n3514), .B2(n3515), .A(net213837), .ZN(net213520) );
  INV_X4 U4980 ( .A(n3517), .ZN(n3514) );
  XNOR2_X2 U4981 ( .A(n3516), .B(n3514), .ZN(net214078) );
  OAI21_X4 U4982 ( .B1(n3518), .B2(n3519), .A(net214083), .ZN(n3517) );
  INV_X4 U4983 ( .A(net214084), .ZN(n3519) );
  INV_X4 U4984 ( .A(net214085), .ZN(n3518) );
  INV_X4 U4985 ( .A(n3515), .ZN(n3516) );
  NAND2_X2 U4986 ( .A1(net214086), .A2(net213837), .ZN(n3515) );
  NAND2_X2 U4987 ( .A1(net214083), .A2(net214085), .ZN(n3520) );
  XNOR2_X2 U4988 ( .A(net214084), .B(n3520), .ZN(net214372) );
  INV_X4 U4989 ( .A(net213818), .ZN(net213514) );
  OAI21_X4 U4990 ( .B1(n3521), .B2(n3522), .A(net213821), .ZN(net213818) );
  INV_X4 U4991 ( .A(net213822), .ZN(n3521) );
  XNOR2_X2 U4992 ( .A(net213822), .B(n3522), .ZN(net214087) );
  NAND2_X4 U4993 ( .A1(net213821), .A2(net214090), .ZN(n3522) );
  OAI211_X2 U4994 ( .C1(n3524), .C2(n3525), .A(net212649), .B(n3425), .ZN(
        net212715) );
  INV_X4 U4995 ( .A(n3523), .ZN(n3525) );
  OAI21_X4 U4996 ( .B1(n3524), .B2(n3525), .A(n3425), .ZN(net213005) );
  OAI21_X4 U4997 ( .B1(n3526), .B2(n3527), .A(net219561), .ZN(n3523) );
  OAI21_X2 U4998 ( .B1(n3526), .B2(n3527), .A(net219561), .ZN(net212656) );
  NAND2_X4 U4999 ( .A1(net213373), .A2(net213374), .ZN(n3528) );
  INV_X2 U5000 ( .A(net213375), .ZN(n3526) );
  OAI21_X2 U5001 ( .B1(net212653), .B2(n3524), .A(n3425), .ZN(net212651) );
  NAND2_X4 U5002 ( .A1(net212700), .A2(n3529), .ZN(net212419) );
  INV_X4 U5003 ( .A(net212704), .ZN(n3531) );
  INV_X4 U5004 ( .A(net212705), .ZN(n3530) );
  NAND2_X2 U5005 ( .A1(n3532), .A2(net214092), .ZN(net214090) );
  NAND2_X2 U5006 ( .A1(a[23]), .A2(net218550), .ZN(n3532) );
  NAND3_X4 U5007 ( .A1(net214093), .A2(a[23]), .A3(net218546), .ZN(net213821)
         );
  INV_X4 U5008 ( .A(net214092), .ZN(net214093) );
  OAI21_X4 U5009 ( .B1(net214101), .B2(n3533), .A(net214103), .ZN(net213822)
         );
  XNOR2_X2 U5010 ( .A(n3533), .B(net214101), .ZN(net220496) );
  NAND2_X4 U5011 ( .A1(net214384), .A2(net214103), .ZN(n3533) );
  OAI21_X4 U5012 ( .B1(n3534), .B2(n3535), .A(net213570), .ZN(net213217) );
  INV_X4 U5013 ( .A(net213571), .ZN(n3535) );
  INV_X1 U5014 ( .A(net213572), .ZN(n3534) );
  XNOR2_X2 U5015 ( .A(net213571), .B(n3536), .ZN(net213740) );
  NOR2_X4 U5016 ( .A1(net241071), .A2(net241074), .ZN(n3537) );
  INV_X4 U5017 ( .A(b[23]), .ZN(net241074) );
  INV_X4 U5018 ( .A(a[6]), .ZN(net241071) );
  XNOR2_X2 U5019 ( .A(n3539), .B(n3540), .ZN(n3538) );
  INV_X4 U5020 ( .A(net212640), .ZN(n3539) );
  INV_X1 U5021 ( .A(n3539), .ZN(net241090) );
  XNOR2_X2 U5022 ( .A(n3540), .B(net212640), .ZN(net241088) );
  NAND2_X2 U5023 ( .A1(b[23]), .A2(a[6]), .ZN(net241082) );
  OAI21_X4 U5024 ( .B1(net213235), .B2(net213236), .A(net213237), .ZN(
        net212930) );
  INV_X4 U5025 ( .A(net213238), .ZN(net213236) );
  INV_X1 U5026 ( .A(net213239), .ZN(net213235) );
  NAND2_X4 U5027 ( .A1(net213237), .A2(net213239), .ZN(net213403) );
  XNOR2_X2 U5028 ( .A(net213403), .B(net213238), .ZN(net213401) );
  NAND2_X4 U5029 ( .A1(net213389), .A2(net213388), .ZN(net213019) );
  INV_X4 U5030 ( .A(net213024), .ZN(net213389) );
  INV_X4 U5031 ( .A(n3541), .ZN(net213024) );
  NAND2_X1 U5032 ( .A1(net213023), .A2(net213024), .ZN(net219749) );
  NAND2_X4 U5033 ( .A1(net213024), .A2(net213023), .ZN(net213384) );
  NAND3_X2 U5034 ( .A1(net213608), .A2(net213609), .A3(n3542), .ZN(net213021)
         );
  NAND2_X2 U5035 ( .A1(net213611), .A2(net213612), .ZN(n3542) );
  INV_X4 U5036 ( .A(net213443), .ZN(net213436) );
  NAND2_X4 U5037 ( .A1(net213751), .A2(net213752), .ZN(net213208) );
  NAND2_X2 U5038 ( .A1(net217552), .A2(net213443), .ZN(net216856) );
  OAI21_X4 U5039 ( .B1(n3543), .B2(n3544), .A(net213532), .ZN(net213115) );
  INV_X4 U5040 ( .A(net213533), .ZN(n3544) );
  INV_X4 U5041 ( .A(net213534), .ZN(n3543) );
  NAND2_X2 U5042 ( .A1(net213532), .A2(net213534), .ZN(n3545) );
  XNOR2_X2 U5043 ( .A(net213533), .B(n3545), .ZN(net213792) );
  OAI21_X4 U5044 ( .B1(n3546), .B2(n3547), .A(net213527), .ZN(net213167) );
  INV_X4 U5045 ( .A(net213528), .ZN(n3547) );
  INV_X4 U5046 ( .A(net213529), .ZN(n3546) );
  XNOR2_X2 U5047 ( .A(net213528), .B(n3548), .ZN(net213797) );
  AOI21_X4 U5048 ( .B1(net213177), .B2(net213178), .A(n3549), .ZN(net213472)
         );
  INV_X4 U5049 ( .A(net213473), .ZN(n3549) );
  XNOR2_X2 U5050 ( .A(net213177), .B(n3550), .ZN(net213782) );
  NAND2_X2 U5051 ( .A1(net213473), .A2(net213178), .ZN(n3550) );
  OAI21_X4 U5052 ( .B1(n3551), .B2(net213541), .A(net213542), .ZN(net213183)
         );
  INV_X2 U5053 ( .A(net213543), .ZN(n3551) );
  INV_X4 U5054 ( .A(net213541), .ZN(net213778) );
  OAI21_X4 U5055 ( .B1(n3552), .B2(net213574), .A(net213575), .ZN(net213222)
         );
  INV_X1 U5056 ( .A(net213579), .ZN(n3552) );
  NAND2_X4 U5057 ( .A1(net213575), .A2(net213579), .ZN(net213737) );
  NAND3_X2 U5058 ( .A1(n3554), .A2(a[23]), .A3(b[4]), .ZN(net213130) );
  XNOR2_X1 U5059 ( .A(net213142), .B(net213140), .ZN(n3554) );
  NAND2_X2 U5060 ( .A1(n3553), .A2(n3555), .ZN(net213132) );
  XOR2_X2 U5061 ( .A(net213142), .B(net213140), .Z(n3555) );
  NAND2_X2 U5062 ( .A1(a[23]), .A2(b[4]), .ZN(n3553) );
  XNOR2_X2 U5063 ( .A(net213804), .B(net213522), .ZN(net213802) );
  INV_X4 U5064 ( .A(net213142), .ZN(net213139) );
  OAI21_X4 U5065 ( .B1(net213139), .B2(net213140), .A(net213141), .ZN(
        net213138) );
  OAI21_X4 U5066 ( .B1(n3557), .B2(n3556), .A(net213546), .ZN(net213190) );
  INV_X2 U5067 ( .A(net213548), .ZN(n3556) );
  INV_X2 U5068 ( .A(n3556), .ZN(n3560) );
  INV_X4 U5069 ( .A(net213547), .ZN(n3557) );
  NAND2_X2 U5070 ( .A1(n3558), .A2(net213775), .ZN(net213191) );
  INV_X4 U5071 ( .A(net213776), .ZN(n3558) );
  NAND2_X4 U5072 ( .A1(net213866), .A2(net213548), .ZN(net214039) );
  NAND2_X2 U5073 ( .A1(net213547), .A2(n3560), .ZN(net213772) );
  NAND2_X2 U5074 ( .A1(n3559), .A2(net213776), .ZN(net213546) );
  OAI21_X4 U5075 ( .B1(net213231), .B2(net213230), .A(net220211), .ZN(
        net212925) );
  INV_X2 U5076 ( .A(net220210), .ZN(net220211) );
  INV_X2 U5077 ( .A(net213232), .ZN(net220210) );
  INV_X2 U5078 ( .A(net213234), .ZN(net213230) );
  INV_X4 U5079 ( .A(net213233), .ZN(net213231) );
  NAND2_X4 U5080 ( .A1(net213232), .A2(net213234), .ZN(net213408) );
  XNOR2_X2 U5081 ( .A(net213233), .B(net213408), .ZN(net213406) );
  NAND2_X2 U5082 ( .A1(n3561), .A2(net213792), .ZN(net213537) );
  INV_X4 U5083 ( .A(net213790), .ZN(n3561) );
  OAI21_X4 U5084 ( .B1(n3562), .B2(n3563), .A(net213850), .ZN(net213538) );
  INV_X4 U5085 ( .A(net213851), .ZN(n3563) );
  INV_X4 U5086 ( .A(net213852), .ZN(n3562) );
  NAND2_X2 U5087 ( .A1(net213790), .A2(net213791), .ZN(net213539) );
  INV_X4 U5088 ( .A(net213792), .ZN(net213791) );
  NAND2_X2 U5089 ( .A1(net213850), .A2(net213852), .ZN(n3564) );
  XNOR2_X2 U5090 ( .A(net213851), .B(n3564), .ZN(net214057) );
  NAND2_X2 U5091 ( .A1(net213513), .A2(n3565), .ZN(net213512) );
  NAND2_X2 U5092 ( .A1(n3566), .A2(net213830), .ZN(n3565) );
  NAND2_X2 U5093 ( .A1(a[25]), .A2(net218558), .ZN(n3566) );
  INV_X4 U5094 ( .A(net213830), .ZN(net217782) );
  AOI21_X4 U5095 ( .B1(net213805), .B2(net213806), .A(n3567), .ZN(net213522)
         );
  INV_X4 U5096 ( .A(net213808), .ZN(n3567) );
  XNOR2_X2 U5097 ( .A(net213805), .B(n3568), .ZN(net214073) );
  NAND2_X2 U5098 ( .A1(net213808), .A2(net213806), .ZN(n3568) );
  NAND3_X2 U5099 ( .A1(net215635), .A2(a[17]), .A3(net218546), .ZN(n5919) );
  XNOR2_X2 U5100 ( .A(net218152), .B(net218153), .ZN(n3569) );
  INV_X1 U5101 ( .A(net214963), .ZN(net223718) );
  XNOR2_X2 U5102 ( .A(n7269), .B(n7127), .ZN(n7130) );
  INV_X2 U5103 ( .A(n7127), .ZN(n7270) );
  OAI21_X2 U5104 ( .B1(net213149), .B2(n7126), .A(n7125), .ZN(n7127) );
  XNOR2_X2 U5105 ( .A(n4908), .B(n4909), .ZN(n3570) );
  NAND2_X2 U5106 ( .A1(n6326), .A2(n6325), .ZN(n6193) );
  INV_X4 U5107 ( .A(n3916), .ZN(n4023) );
  NAND2_X2 U5108 ( .A1(n3342), .A2(net216840), .ZN(n4884) );
  INV_X2 U5109 ( .A(n3867), .ZN(n3865) );
  INV_X2 U5110 ( .A(n6325), .ZN(n6329) );
  NAND2_X4 U5111 ( .A1(n3966), .A2(n5942), .ZN(n5949) );
  NAND2_X4 U5112 ( .A1(n6027), .A2(n6153), .ZN(n6072) );
  OAI21_X2 U5113 ( .B1(net217288), .B2(net217287), .A(net219864), .ZN(
        net217106) );
  NAND3_X2 U5114 ( .A1(net214571), .A2(net220181), .A3(net214570), .ZN(
        net214568) );
  NAND2_X4 U5115 ( .A1(net218556), .A2(a[5]), .ZN(n4051) );
  NAND2_X1 U5116 ( .A1(net224032), .A2(net218116), .ZN(n4098) );
  INV_X2 U5117 ( .A(n4093), .ZN(n4065) );
  NAND2_X4 U5118 ( .A1(n4102), .A2(n4101), .ZN(n4096) );
  NAND2_X4 U5119 ( .A1(n4035), .A2(n4034), .ZN(net218272) );
  INV_X8 U5120 ( .A(net218238), .ZN(net223234) );
  INV_X2 U5121 ( .A(net241371), .ZN(net241372) );
  NAND2_X4 U5122 ( .A1(net241364), .A2(net241365), .ZN(n3573) );
  NAND2_X4 U5123 ( .A1(net241366), .A2(n3573), .ZN(net218156) );
  INV_X4 U5124 ( .A(net218158), .ZN(net241364) );
  NAND2_X4 U5125 ( .A1(net218157), .A2(net218156), .ZN(net218095) );
  NAND2_X2 U5126 ( .A1(n6833), .A2(n6832), .ZN(n3574) );
  NAND2_X2 U5127 ( .A1(n3575), .A2(n6962), .ZN(n6839) );
  INV_X4 U5128 ( .A(n3574), .ZN(n3575) );
  NAND2_X2 U5129 ( .A1(n6830), .A2(n6829), .ZN(n3578) );
  NAND2_X4 U5130 ( .A1(n3576), .A2(n3577), .ZN(n3579) );
  NAND2_X4 U5131 ( .A1(n3578), .A2(n3579), .ZN(n6831) );
  INV_X4 U5132 ( .A(n6830), .ZN(n3576) );
  INV_X4 U5133 ( .A(n6829), .ZN(n3577) );
  NAND2_X4 U5134 ( .A1(n3580), .A2(n3581), .ZN(n3583) );
  INV_X4 U5135 ( .A(net215064), .ZN(n3580) );
  INV_X4 U5136 ( .A(n6085), .ZN(n3581) );
  INV_X2 U5137 ( .A(n6839), .ZN(n6834) );
  NAND2_X4 U5138 ( .A1(n6953), .A2(n6831), .ZN(n6838) );
  INV_X2 U5139 ( .A(n4736), .ZN(n4740) );
  NAND2_X4 U5140 ( .A1(n4737), .A2(n4736), .ZN(n4738) );
  INV_X4 U5141 ( .A(net218337), .ZN(net217879) );
  INV_X8 U5142 ( .A(net215428), .ZN(net215426) );
  OAI21_X4 U5143 ( .B1(n3739), .B2(n3741), .A(n3738), .ZN(n3740) );
  NAND2_X2 U5144 ( .A1(n3814), .A2(n3813), .ZN(n5206) );
  INV_X2 U5145 ( .A(n4981), .ZN(n4985) );
  XNOR2_X2 U5146 ( .A(net214603), .B(n3805), .ZN(n6384) );
  NOR2_X2 U5147 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  INV_X4 U5148 ( .A(n5087), .ZN(n4980) );
  INV_X8 U5149 ( .A(n3618), .ZN(n3615) );
  NAND2_X4 U5150 ( .A1(n3924), .A2(n6825), .ZN(net213612) );
  NAND2_X2 U5151 ( .A1(n3584), .A2(net217233), .ZN(n3586) );
  NAND2_X2 U5152 ( .A1(n3585), .A2(n3586), .ZN(n4127) );
  INV_X2 U5153 ( .A(net218054), .ZN(n3584) );
  OAI21_X2 U5154 ( .B1(n5770), .B2(n5769), .A(net215477), .ZN(net215675) );
  CLKBUF_X3 U5155 ( .A(n3615), .Z(n3587) );
  NAND2_X4 U5156 ( .A1(net217072), .A2(net217071), .ZN(net216839) );
  NAND3_X2 U5157 ( .A1(net219934), .A2(net215516), .A3(net215517), .ZN(n5980)
         );
  INV_X2 U5158 ( .A(net214710), .ZN(n3588) );
  CLKBUF_X3 U5159 ( .A(n6148), .Z(n3941) );
  INV_X2 U5160 ( .A(net219178), .ZN(net214457) );
  NAND2_X2 U5161 ( .A1(n3589), .A2(n3590), .ZN(n3592) );
  NAND2_X2 U5162 ( .A1(n3591), .A2(n3592), .ZN(n6221) );
  INV_X4 U5163 ( .A(n6383), .ZN(n3589) );
  NAND2_X4 U5164 ( .A1(b[11]), .A2(a[11]), .ZN(n6382) );
  INV_X2 U5165 ( .A(net215477), .ZN(n3721) );
  INV_X2 U5166 ( .A(n6838), .ZN(n6835) );
  OAI21_X2 U5167 ( .B1(n6087), .B2(n6088), .A(n6428), .ZN(n6092) );
  NAND2_X4 U5168 ( .A1(n6308), .A2(n6152), .ZN(n6077) );
  NAND2_X4 U5169 ( .A1(n6061), .A2(n6062), .ZN(n6159) );
  NAND2_X4 U5170 ( .A1(n5656), .A2(net215848), .ZN(n5785) );
  NAND3_X4 U5171 ( .A1(n6039), .A2(a[18]), .A3(net218536), .ZN(n6335) );
  NAND2_X2 U5172 ( .A1(net215218), .A2(net215219), .ZN(net214857) );
  INV_X8 U5173 ( .A(n4729), .ZN(n4733) );
  XNOR2_X2 U5174 ( .A(n4932), .B(n3594), .ZN(n3593) );
  AND3_X4 U5175 ( .A1(n4966), .A2(n4965), .A3(n4964), .ZN(n3594) );
  INV_X4 U5176 ( .A(n6701), .ZN(n6702) );
  NAND2_X4 U5177 ( .A1(net213743), .A2(n6932), .ZN(net213572) );
  OAI21_X4 U5178 ( .B1(net213766), .B2(n6714), .A(net213553), .ZN(n6781) );
  XNOR2_X2 U5179 ( .A(n5828), .B(n5831), .ZN(n3595) );
  OAI21_X2 U5180 ( .B1(n6019), .B2(n6018), .A(net215224), .ZN(net214972) );
  NAND2_X4 U5181 ( .A1(n6505), .A2(n6504), .ZN(n6786) );
  NAND2_X4 U5182 ( .A1(n4902), .A2(n4901), .ZN(n5092) );
  NAND2_X4 U5183 ( .A1(n5349), .A2(n5348), .ZN(n5522) );
  INV_X4 U5184 ( .A(n5471), .ZN(n5345) );
  AOI21_X4 U5185 ( .B1(net216392), .B2(net216219), .A(net216221), .ZN(
        net216400) );
  INV_X4 U5186 ( .A(net216653), .ZN(net216649) );
  NAND2_X2 U5187 ( .A1(n5635), .A2(n5636), .ZN(n5910) );
  NAND2_X4 U5188 ( .A1(n6754), .A2(n6753), .ZN(n6911) );
  NAND2_X4 U5189 ( .A1(net214059), .A2(n6760), .ZN(n6906) );
  NAND2_X4 U5190 ( .A1(n5819), .A2(n5820), .ZN(net215335) );
  INV_X4 U5191 ( .A(n3424), .ZN(n6248) );
  INV_X2 U5192 ( .A(n5664), .ZN(n3908) );
  NAND2_X4 U5193 ( .A1(n5948), .A2(n5943), .ZN(n5674) );
  NAND2_X4 U5194 ( .A1(n5348), .A2(n5521), .ZN(n5129) );
  OAI21_X4 U5195 ( .B1(net220385), .B2(net215206), .A(net215199), .ZN(n3732)
         );
  NAND2_X4 U5196 ( .A1(n3691), .A2(net216576), .ZN(net216583) );
  OAI21_X4 U5197 ( .B1(net219339), .B2(net216657), .A(net216658), .ZN(n3691)
         );
  INV_X4 U5198 ( .A(net223819), .ZN(net218215) );
  NAND2_X4 U5199 ( .A1(n5401), .A2(n5400), .ZN(n5472) );
  INV_X8 U5200 ( .A(net220396), .ZN(net218334) );
  NAND2_X2 U5201 ( .A1(net216759), .A2(net216760), .ZN(n3599) );
  NAND2_X4 U5202 ( .A1(n3597), .A2(n3598), .ZN(n3600) );
  NAND2_X4 U5203 ( .A1(n3600), .A2(n3599), .ZN(n5006) );
  INV_X8 U5204 ( .A(net216759), .ZN(n3597) );
  INV_X4 U5205 ( .A(net216760), .ZN(n3598) );
  INV_X2 U5206 ( .A(n5006), .ZN(n5003) );
  NAND2_X4 U5207 ( .A1(n4061), .A2(n4060), .ZN(n4062) );
  INV_X4 U5208 ( .A(n5433), .ZN(n5431) );
  INV_X4 U5209 ( .A(n5207), .ZN(n5071) );
  NAND2_X2 U5210 ( .A1(n4147), .A2(n4152), .ZN(n4148) );
  NAND2_X4 U5211 ( .A1(n6743), .A2(n6548), .ZN(n6744) );
  XNOR2_X1 U5212 ( .A(n5384), .B(n5383), .ZN(n3964) );
  NAND3_X4 U5213 ( .A1(a[22]), .A2(net214385), .A3(net218548), .ZN(net214103)
         );
  OAI21_X2 U5214 ( .B1(net214726), .B2(net219162), .A(net214727), .ZN(
        net214723) );
  NAND2_X4 U5215 ( .A1(n7015), .A2(net213508), .ZN(n7114) );
  NAND2_X4 U5216 ( .A1(n7253), .A2(n7254), .ZN(n7161) );
  NAND2_X4 U5217 ( .A1(n7260), .A2(n7259), .ZN(n7152) );
  OAI21_X4 U5218 ( .B1(n3676), .B2(n3677), .A(net215445), .ZN(n3683) );
  INV_X8 U5219 ( .A(net215330), .ZN(n3664) );
  NAND2_X4 U5220 ( .A1(net214960), .A2(net214961), .ZN(net215354) );
  NAND2_X4 U5221 ( .A1(n3729), .A2(n3728), .ZN(net214961) );
  NAND2_X4 U5222 ( .A1(n6076), .A2(n6075), .ZN(n6152) );
  NAND2_X4 U5223 ( .A1(n5662), .A2(n5780), .ZN(n5777) );
  NAND3_X4 U5224 ( .A1(n5661), .A2(a[15]), .A3(net218534), .ZN(n5780) );
  NOR2_X4 U5225 ( .A1(n3662), .A2(n3602), .ZN(n3601) );
  NOR2_X4 U5226 ( .A1(n3694), .A2(n3695), .ZN(n3692) );
  INV_X4 U5227 ( .A(n3771), .ZN(n6803) );
  NAND2_X4 U5228 ( .A1(net215334), .A2(net215335), .ZN(net215338) );
  INV_X4 U5229 ( .A(n5558), .ZN(n5560) );
  INV_X4 U5230 ( .A(n4094), .ZN(n4102) );
  INV_X8 U5231 ( .A(n4011), .ZN(n4033) );
  NAND2_X2 U5232 ( .A1(n6490), .A2(n6489), .ZN(n6688) );
  NAND2_X1 U5233 ( .A1(n6694), .A2(n6693), .ZN(n6696) );
  INV_X2 U5234 ( .A(net215334), .ZN(n3665) );
  INV_X2 U5235 ( .A(n5772), .ZN(n3604) );
  INV_X4 U5236 ( .A(n3604), .ZN(n3605) );
  INV_X4 U5237 ( .A(n5215), .ZN(n5217) );
  INV_X4 U5238 ( .A(n6588), .ZN(n6586) );
  NAND2_X4 U5239 ( .A1(n5814), .A2(n5815), .ZN(n5962) );
  NAND2_X4 U5240 ( .A1(net216210), .A2(net219220), .ZN(n3861) );
  NAND2_X2 U5241 ( .A1(n5474), .A2(n5638), .ZN(n5393) );
  NAND2_X4 U5242 ( .A1(b[1]), .A2(a[1]), .ZN(n3606) );
  INV_X4 U5243 ( .A(n4029), .ZN(n4071) );
  NAND2_X4 U5244 ( .A1(n4007), .A2(n4029), .ZN(n4046) );
  INV_X1 U5245 ( .A(net215583), .ZN(net215780) );
  INV_X8 U5246 ( .A(net213729), .ZN(net213724) );
  INV_X8 U5247 ( .A(n5614), .ZN(n3932) );
  NAND2_X2 U5248 ( .A1(n3815), .A2(n5209), .ZN(n5131) );
  NAND2_X4 U5249 ( .A1(n3855), .A2(n3854), .ZN(n3845) );
  INV_X2 U5250 ( .A(net214434), .ZN(n3851) );
  NAND2_X4 U5251 ( .A1(n6795), .A2(n6794), .ZN(n6892) );
  INV_X4 U5252 ( .A(net212645), .ZN(net241055) );
  NOR2_X2 U5253 ( .A1(net241076), .A2(net241077), .ZN(net212452) );
  NAND2_X4 U5254 ( .A1(n3607), .A2(net214958), .ZN(net215353) );
  XNOR2_X2 U5255 ( .A(net215353), .B(net215354), .ZN(net215350) );
  AOI21_X2 U5256 ( .B1(net215353), .B2(net214960), .A(net214954), .ZN(
        net215129) );
  OAI21_X4 U5257 ( .B1(net215426), .B2(net215425), .A(net215427), .ZN(n3607)
         );
  INV_X2 U5258 ( .A(net215429), .ZN(net215425) );
  OAI21_X2 U5259 ( .B1(net215426), .B2(net215425), .A(net215427), .ZN(
        net223455) );
  INV_X2 U5260 ( .A(net215425), .ZN(net219611) );
  OAI21_X4 U5261 ( .B1(net215665), .B2(net215664), .A(net215666), .ZN(
        net215428) );
  INV_X8 U5262 ( .A(net215587), .ZN(net215666) );
  OAI21_X2 U5263 ( .B1(net215665), .B2(net215664), .A(net215666), .ZN(
        net223706) );
  INV_X1 U5264 ( .A(net215669), .ZN(net215664) );
  NAND2_X4 U5265 ( .A1(net215431), .A2(net215430), .ZN(net214958) );
  NAND2_X4 U5266 ( .A1(net215427), .A2(net214958), .ZN(net215593) );
  INV_X4 U5267 ( .A(net215595), .ZN(net215430) );
  NAND2_X4 U5268 ( .A1(n3608), .A2(net215595), .ZN(net215427) );
  NAND2_X4 U5269 ( .A1(n3613), .A2(n3609), .ZN(net215429) );
  NAND2_X1 U5270 ( .A1(net215429), .A2(net215667), .ZN(net215798) );
  NAND2_X4 U5271 ( .A1(net215667), .A2(net215429), .ZN(net215587) );
  INV_X4 U5272 ( .A(net215802), .ZN(n3609) );
  XNOR2_X2 U5273 ( .A(net215805), .B(n3610), .ZN(n3613) );
  NOR2_X4 U5274 ( .A1(n3611), .A2(n3612), .ZN(n3610) );
  NOR2_X4 U5275 ( .A1(n3611), .A2(n3612), .ZN(net219656) );
  INV_X4 U5276 ( .A(net215363), .ZN(n3611) );
  NAND2_X1 U5277 ( .A1(net215587), .A2(net215799), .ZN(net223270) );
  NOR2_X4 U5278 ( .A1(net218277), .A2(n3615), .ZN(n3614) );
  OAI21_X4 U5279 ( .B1(n3614), .B2(net220033), .A(net218272), .ZN(net218270)
         );
  AOI21_X2 U5280 ( .B1(n3615), .B2(net218276), .A(net218277), .ZN(net218308)
         );
  NAND2_X4 U5281 ( .A1(net217879), .A2(n3305), .ZN(n3618) );
  MUX2_X2 U5282 ( .A(net217877), .B(net217878), .S(net217879), .Z(net217876)
         );
  XNOR2_X2 U5283 ( .A(n3619), .B(net218339), .ZN(net218337) );
  NAND2_X2 U5284 ( .A1(a[0]), .A2(a[1]), .ZN(n3620) );
  XNOR2_X2 U5285 ( .A(net217857), .B(n3606), .ZN(n3619) );
  AND2_X2 U5286 ( .A1(net217857), .A2(net218354), .ZN(net218362) );
  INV_X4 U5287 ( .A(net218297), .ZN(net218277) );
  INV_X4 U5288 ( .A(net218277), .ZN(net220153) );
  NAND3_X2 U5289 ( .A1(net218322), .A2(net218321), .A3(n3616), .ZN(net218297)
         );
  INV_X2 U5290 ( .A(n3617), .ZN(n3616) );
  AOI21_X4 U5291 ( .B1(net218322), .B2(net218321), .A(n3616), .ZN(net220033)
         );
  NAND2_X1 U5292 ( .A1(net218550), .A2(net218480), .ZN(n3617) );
  OAI22_X4 U5293 ( .A1(net220395), .A2(net220394), .B1(net220395), .B2(
        net218367), .ZN(net218352) );
  NOR2_X4 U5294 ( .A1(net214819), .A2(n3621), .ZN(n3622) );
  AOI21_X4 U5295 ( .B1(n3622), .B2(net214817), .A(net214717), .ZN(net214815)
         );
  INV_X4 U5296 ( .A(net214820), .ZN(n3621) );
  AOI21_X4 U5297 ( .B1(net214720), .B2(net214721), .A(n3621), .ZN(net214718)
         );
  INV_X2 U5298 ( .A(n3621), .ZN(net219530) );
  NAND2_X2 U5299 ( .A1(n3623), .A2(net215300), .ZN(net214820) );
  NAND2_X4 U5300 ( .A1(net214721), .A2(net214820), .ZN(net215298) );
  INV_X4 U5301 ( .A(net215301), .ZN(n3623) );
  OAI21_X2 U5302 ( .B1(net214717), .B2(net214718), .A(net214719), .ZN(
        net214715) );
  INV_X4 U5303 ( .A(net215076), .ZN(net215074) );
  INV_X4 U5304 ( .A(net215300), .ZN(net215302) );
  NAND2_X4 U5305 ( .A1(net215302), .A2(net215301), .ZN(net214721) );
  NAND2_X4 U5306 ( .A1(net215077), .A2(net215076), .ZN(net214818) );
  NAND2_X2 U5307 ( .A1(b[22]), .A2(a[5]), .ZN(net213388) );
  INV_X2 U5308 ( .A(net213388), .ZN(net213023) );
  XNOR2_X2 U5309 ( .A(net213397), .B(net213398), .ZN(net220449) );
  INV_X4 U5310 ( .A(net213394), .ZN(net213396) );
  NAND2_X4 U5311 ( .A1(net213393), .A2(net213394), .ZN(net213033) );
  INV_X4 U5312 ( .A(net213395), .ZN(net213393) );
  XNOR2_X2 U5313 ( .A(net213397), .B(net213398), .ZN(net213395) );
  AOI21_X4 U5314 ( .B1(net213604), .B2(net213605), .A(net213606), .ZN(
        net213031) );
  INV_X4 U5315 ( .A(net213607), .ZN(net213606) );
  NAND2_X2 U5316 ( .A1(a[5]), .A2(b[21]), .ZN(net213603) );
  NAND2_X4 U5317 ( .A1(net218103), .A2(net217107), .ZN(net218104) );
  AOI22_X2 U5318 ( .A1(net218101), .A2(net219864), .B1(net218104), .B2(
        net218103), .ZN(net218071) );
  XNOR2_X2 U5319 ( .A(net218110), .B(n3174), .ZN(net217246) );
  CLKBUF_X3 U5320 ( .A(net217107), .Z(net219368) );
  NAND2_X2 U5321 ( .A1(net217107), .A2(net218105), .ZN(net218149) );
  NAND2_X4 U5322 ( .A1(net218112), .A2(net218111), .ZN(net218103) );
  INV_X4 U5323 ( .A(net218151), .ZN(net218111) );
  NAND2_X4 U5324 ( .A1(net218112), .A2(net218111), .ZN(net218105) );
  INV_X4 U5325 ( .A(net218150), .ZN(net218112) );
  NAND2_X4 U5326 ( .A1(net214587), .A2(net214970), .ZN(net215097) );
  XNOR2_X2 U5327 ( .A(net215097), .B(net215096), .ZN(net215093) );
  XNOR2_X2 U5328 ( .A(net215097), .B(net215096), .ZN(net223508) );
  NAND2_X4 U5329 ( .A1(net215101), .A2(net215100), .ZN(net214587) );
  NAND2_X2 U5330 ( .A1(net214588), .A2(net214587), .ZN(net214846) );
  NAND2_X2 U5331 ( .A1(net214586), .A2(net214587), .ZN(net214584) );
  INV_X2 U5332 ( .A(net215099), .ZN(net215101) );
  NAND2_X2 U5333 ( .A1(net215098), .A2(net215099), .ZN(net214970) );
  NAND3_X2 U5334 ( .A1(net214970), .A2(net223712), .A3(net214972), .ZN(
        net214588) );
  INV_X4 U5335 ( .A(net215100), .ZN(net215098) );
  NAND2_X2 U5336 ( .A1(net214878), .A2(net215123), .ZN(net215348) );
  NAND2_X4 U5337 ( .A1(net215352), .A2(net215351), .ZN(net214878) );
  NAND2_X1 U5338 ( .A1(net214878), .A2(net223182), .ZN(net215212) );
  INV_X4 U5339 ( .A(net215350), .ZN(net215352) );
  NAND2_X2 U5340 ( .A1(net215350), .A2(net215349), .ZN(net215123) );
  INV_X4 U5341 ( .A(net215123), .ZN(net214879) );
  INV_X4 U5342 ( .A(net215351), .ZN(net215349) );
  NAND2_X4 U5343 ( .A1(net214975), .A2(net214714), .ZN(net215091) );
  XNOR2_X2 U5344 ( .A(net215091), .B(net215088), .ZN(net223874) );
  NAND2_X4 U5345 ( .A1(net215095), .A2(net215094), .ZN(net214975) );
  OAI21_X4 U5346 ( .B1(net214973), .B2(net214974), .A(net214975), .ZN(
        net214713) );
  INV_X4 U5347 ( .A(net215093), .ZN(net215095) );
  NAND2_X4 U5348 ( .A1(net215092), .A2(net223508), .ZN(net214714) );
  INV_X4 U5349 ( .A(net215094), .ZN(net215092) );
  NAND2_X2 U5350 ( .A1(a[6]), .A2(b[21]), .ZN(net213394) );
  NAND2_X4 U5351 ( .A1(net213595), .A2(net220046), .ZN(net213397) );
  INV_X4 U5352 ( .A(net218066), .ZN(net218065) );
  NAND2_X2 U5353 ( .A1(net218068), .A2(net218067), .ZN(net216946) );
  INV_X2 U5354 ( .A(net218069), .ZN(net218068) );
  NAND2_X2 U5355 ( .A1(net218067), .A2(net218068), .ZN(net223932) );
  INV_X4 U5356 ( .A(net218070), .ZN(net218067) );
  NAND2_X2 U5357 ( .A1(net218070), .A2(net218069), .ZN(net217243) );
  NAND2_X4 U5358 ( .A1(net218809), .A2(net217243), .ZN(net216944) );
  XNOR2_X2 U5359 ( .A(net218071), .B(net218072), .ZN(net218069) );
  NAND2_X2 U5360 ( .A1(b[4]), .A2(a[5]), .ZN(net218070) );
  INV_X32 U5361 ( .A(a[5]), .ZN(net218456) );
  NAND2_X4 U5362 ( .A1(net218101), .A2(net218106), .ZN(net218110) );
  NAND2_X2 U5363 ( .A1(net218538), .A2(a[5]), .ZN(net218151) );
  XNOR2_X2 U5364 ( .A(net218152), .B(net218153), .ZN(net218150) );
  NAND2_X2 U5365 ( .A1(net217262), .A2(net218095), .ZN(net218153) );
  OAI22_X4 U5366 ( .A1(net218170), .A2(net218099), .B1(net218172), .B2(
        net218171), .ZN(net218152) );
  INV_X4 U5367 ( .A(net218098), .ZN(net218171) );
  AOI21_X4 U5368 ( .B1(net218173), .B2(net218174), .A(net218175), .ZN(
        net218172) );
  INV_X8 U5369 ( .A(net218100), .ZN(net218175) );
  INV_X2 U5370 ( .A(net218175), .ZN(net219065) );
  NAND2_X2 U5371 ( .A1(net217261), .A2(net217262), .ZN(net218093) );
  NAND2_X4 U5372 ( .A1(net218095), .A2(net218094), .ZN(net217261) );
  OAI211_X4 U5373 ( .C1(net218170), .C2(net217258), .A(net217259), .B(
        net217260), .ZN(net217118) );
  XNOR2_X2 U5374 ( .A(net218268), .B(net218239), .ZN(net218234) );
  XNOR2_X2 U5375 ( .A(net218238), .B(net218239), .ZN(net218237) );
  NAND2_X4 U5376 ( .A1(net223819), .A2(net218098), .ZN(net218170) );
  NAND2_X2 U5377 ( .A1(net213402), .A2(net213401), .ZN(net213242) );
  INV_X4 U5378 ( .A(net213400), .ZN(net213402) );
  NAND2_X4 U5379 ( .A1(net213399), .A2(net213400), .ZN(net213248) );
  INV_X4 U5380 ( .A(net213401), .ZN(net213399) );
  NAND2_X2 U5381 ( .A1(n3624), .A2(net214855), .ZN(net215103) );
  XNOR2_X2 U5382 ( .A(net215103), .B(net215102), .ZN(net215099) );
  NAND2_X2 U5383 ( .A1(net215107), .A2(net215106), .ZN(net223422) );
  NAND2_X2 U5384 ( .A1(net215104), .A2(net215105), .ZN(net214855) );
  NAND3_X2 U5385 ( .A1(net214855), .A2(net214856), .A3(net214857), .ZN(
        net214853) );
  INV_X4 U5386 ( .A(net215106), .ZN(net215104) );
  NAND2_X2 U5387 ( .A1(b[12]), .A2(a[9]), .ZN(net215106) );
  XNOR2_X2 U5388 ( .A(n3625), .B(n3626), .ZN(net215105) );
  NAND2_X2 U5389 ( .A1(net214864), .A2(net214968), .ZN(n3626) );
  NAND2_X4 U5390 ( .A1(net215213), .A2(net220004), .ZN(n3625) );
  CLKBUF_X3 U5391 ( .A(net214969), .Z(net220004) );
  INV_X2 U5392 ( .A(net214967), .ZN(net215213) );
  INV_X2 U5393 ( .A(net214864), .ZN(net219770) );
  OAI21_X2 U5394 ( .B1(net214966), .B2(net214967), .A(net214968), .ZN(
        net214863) );
  INV_X1 U5395 ( .A(net214969), .ZN(net214966) );
  NAND2_X4 U5396 ( .A1(net214797), .A2(net214796), .ZN(net214543) );
  NAND2_X4 U5397 ( .A1(net214543), .A2(net214542), .ZN(net214793) );
  INV_X2 U5398 ( .A(net214795), .ZN(net214797) );
  NAND2_X2 U5399 ( .A1(b[18]), .A2(net219055), .ZN(net214796) );
  INV_X4 U5400 ( .A(net214796), .ZN(net214794) );
  INV_X32 U5401 ( .A(net219069), .ZN(net219055) );
  INV_X32 U5402 ( .A(a[4]), .ZN(net219069) );
  XNOR2_X2 U5403 ( .A(net217990), .B(net219069), .ZN(net217761) );
  NAND2_X2 U5404 ( .A1(net214794), .A2(net214795), .ZN(net214542) );
  NOR2_X4 U5405 ( .A1(net214808), .A2(net214809), .ZN(n3627) );
  INV_X4 U5406 ( .A(net214724), .ZN(net214809) );
  AOI21_X2 U5407 ( .B1(n3629), .B2(n3630), .A(n3631), .ZN(n3628) );
  INV_X4 U5408 ( .A(net214727), .ZN(n3631) );
  NOR2_X4 U5409 ( .A1(n3631), .A2(net219162), .ZN(net215064) );
  NOR2_X2 U5410 ( .A1(n3633), .A2(n3634), .ZN(n3632) );
  INV_X4 U5411 ( .A(net214731), .ZN(n3634) );
  INV_X4 U5412 ( .A(net214732), .ZN(n3633) );
  INV_X1 U5413 ( .A(n3633), .ZN(net219934) );
  OAI21_X4 U5414 ( .B1(net215519), .B2(n3633), .A(net215518), .ZN(net215282)
         );
  INV_X2 U5415 ( .A(net224078), .ZN(n3635) );
  NAND2_X4 U5416 ( .A1(b[0]), .A2(a[4]), .ZN(net219063) );
  NAND2_X2 U5417 ( .A1(net214723), .A2(net214724), .ZN(net214460) );
  NAND2_X4 U5418 ( .A1(net214460), .A2(net214461), .ZN(net214551) );
  NAND2_X4 U5419 ( .A1(net219429), .A2(net214812), .ZN(net214461) );
  INV_X4 U5420 ( .A(net214811), .ZN(net214812) );
  NAND2_X2 U5421 ( .A1(b[17]), .A2(a[5]), .ZN(net214811) );
  NAND2_X4 U5422 ( .A1(net214810), .A2(net214811), .ZN(net214724) );
  NOR2_X4 U5423 ( .A1(n3636), .A2(net219178), .ZN(net214814) );
  XNOR2_X2 U5424 ( .A(net214815), .B(net214814), .ZN(net214810) );
  INV_X4 U5425 ( .A(net214716), .ZN(n3636) );
  NAND2_X4 U5426 ( .A1(net214715), .A2(net214716), .ZN(net214456) );
  NAND2_X4 U5427 ( .A1(net214817), .A2(net219530), .ZN(net215072) );
  NAND2_X4 U5428 ( .A1(b[0]), .A2(a[2]), .ZN(net217790) );
  MUX2_X2 U5429 ( .A(net219063), .B(n3881), .S(net218558), .Z(net217972) );
  NAND2_X4 U5430 ( .A1(n3637), .A2(n3322), .ZN(net215669) );
  NAND2_X2 U5431 ( .A1(net215668), .A2(n3281), .ZN(net215586) );
  OAI21_X4 U5432 ( .B1(n3322), .B2(net219336), .A(net215669), .ZN(net215796)
         );
  NAND2_X2 U5433 ( .A1(net215814), .A2(net215809), .ZN(net216016) );
  XNOR2_X1 U5434 ( .A(net216016), .B(net216017), .ZN(net219336) );
  NAND3_X4 U5435 ( .A1(net215807), .A2(n3638), .A3(net215812), .ZN(net216017)
         );
  INV_X4 U5436 ( .A(net215810), .ZN(n3638) );
  INV_X2 U5437 ( .A(net215813), .ZN(net215810) );
  NOR2_X4 U5438 ( .A1(net215811), .A2(net215810), .ZN(net215806) );
  INV_X2 U5439 ( .A(net215814), .ZN(net215661) );
  INV_X4 U5440 ( .A(net215809), .ZN(net215808) );
  AOI21_X4 U5441 ( .B1(net215806), .B2(net215807), .A(net215808), .ZN(
        net215662) );
  NAND2_X2 U5442 ( .A1(b[14]), .A2(a[7]), .ZN(net215094) );
  NAND2_X4 U5443 ( .A1(net214971), .A2(net215224), .ZN(net215316) );
  CLKBUF_X2 U5444 ( .A(net214971), .Z(net223712) );
  NAND2_X4 U5445 ( .A1(net215084), .A2(net215083), .ZN(net214570) );
  NAND2_X4 U5446 ( .A1(n3639), .A2(net214570), .ZN(net215082) );
  INV_X4 U5447 ( .A(net215085), .ZN(net215083) );
  XNOR2_X2 U5448 ( .A(net215087), .B(net215088), .ZN(net215084) );
  NAND2_X2 U5449 ( .A1(b[15]), .A2(a[6]), .ZN(net215085) );
  AOI21_X4 U5450 ( .B1(net215089), .B2(net214979), .A(net214973), .ZN(
        net215088) );
  INV_X4 U5451 ( .A(net215090), .ZN(net214973) );
  XNOR2_X2 U5452 ( .A(net215089), .B(net215310), .ZN(net223908) );
  INV_X4 U5453 ( .A(net214979), .ZN(net214978) );
  NAND2_X2 U5454 ( .A1(net214979), .A2(net215090), .ZN(net215310) );
  NAND2_X2 U5455 ( .A1(b[13]), .A2(a[8]), .ZN(net215100) );
  NAND2_X2 U5456 ( .A1(net214856), .A2(net214857), .ZN(net215102) );
  NAND2_X4 U5457 ( .A1(net215219), .A2(net214856), .ZN(net215322) );
  NAND2_X2 U5458 ( .A1(net214179), .A2(net214178), .ZN(net214175) );
  AOI21_X4 U5459 ( .B1(net214175), .B2(net214174), .A(n3601), .ZN(net213891)
         );
  OAI21_X4 U5460 ( .B1(n3641), .B2(net214541), .A(net214542), .ZN(net214179)
         );
  AOI21_X2 U5461 ( .B1(net214179), .B2(net214178), .A(net220149), .ZN(
        net214289) );
  XNOR2_X2 U5462 ( .A(net214179), .B(net214539), .ZN(net214536) );
  INV_X4 U5463 ( .A(n3642), .ZN(n3641) );
  NAND2_X4 U5464 ( .A1(net214545), .A2(net214546), .ZN(n3642) );
  NAND2_X2 U5465 ( .A1(n3644), .A2(net214549), .ZN(net214178) );
  NAND2_X4 U5466 ( .A1(net214178), .A2(net214174), .ZN(net214539) );
  INV_X4 U5467 ( .A(n3643), .ZN(n3644) );
  NOR2_X4 U5468 ( .A1(n3644), .A2(net214549), .ZN(net220149) );
  XNOR2_X2 U5469 ( .A(n3645), .B(net214551), .ZN(n3643) );
  NAND2_X4 U5470 ( .A1(net213992), .A2(net214459), .ZN(n3645) );
  NAND2_X4 U5471 ( .A1(net214786), .A2(net214545), .ZN(net215059) );
  NAND2_X1 U5472 ( .A1(net214786), .A2(net214545), .ZN(net214784) );
  NAND2_X2 U5473 ( .A1(net214546), .A2(net214545), .ZN(net214792) );
  NAND2_X4 U5474 ( .A1(n3640), .A2(net213992), .ZN(net213989) );
  OAI21_X4 U5475 ( .B1(net216768), .B2(net219256), .A(net216831), .ZN(
        net216777) );
  XNOR2_X2 U5476 ( .A(net216777), .B(net216282), .ZN(net216775) );
  OAI21_X2 U5477 ( .B1(net216832), .B2(net216833), .A(net216834), .ZN(
        net216831) );
  NOR2_X4 U5478 ( .A1(net216830), .A2(net216770), .ZN(net216834) );
  INV_X8 U5479 ( .A(net216646), .ZN(net216770) );
  AOI21_X4 U5480 ( .B1(net216771), .B2(net216651), .A(net216770), .ZN(
        net216978) );
  NOR2_X1 U5481 ( .A1(net216770), .A2(net216771), .ZN(net216769) );
  INV_X4 U5482 ( .A(net216648), .ZN(net216830) );
  INV_X2 U5483 ( .A(net216771), .ZN(net216833) );
  INV_X2 U5484 ( .A(net216651), .ZN(net216832) );
  INV_X2 U5485 ( .A(net219713), .ZN(net219256) );
  INV_X4 U5486 ( .A(net216835), .ZN(net216768) );
  NAND2_X4 U5487 ( .A1(n3648), .A2(n3647), .ZN(net216646) );
  NAND2_X2 U5488 ( .A1(net216651), .A2(net216646), .ZN(net217078) );
  OAI221_X4 U5489 ( .B1(n3649), .B2(net216646), .C1(net216645), .C2(net216647), 
        .A(net219713), .ZN(net216285) );
  INV_X4 U5490 ( .A(net217088), .ZN(n3647) );
  XOR2_X2 U5491 ( .A(net217092), .B(net217091), .Z(n3648) );
  NAND2_X4 U5492 ( .A1(net216936), .A2(n3646), .ZN(net216648) );
  NAND2_X2 U5493 ( .A1(net216648), .A2(net219641), .ZN(net216835) );
  INV_X4 U5494 ( .A(net216934), .ZN(n3646) );
  NAND2_X2 U5495 ( .A1(n3646), .A2(net216936), .ZN(net219713) );
  NAND2_X4 U5496 ( .A1(net217079), .A2(net216652), .ZN(net216771) );
  XNOR2_X2 U5497 ( .A(net217078), .B(net216771), .ZN(net217075) );
  NAND3_X2 U5498 ( .A1(net217086), .A2(net219494), .A3(net217084), .ZN(
        net217079) );
  INV_X4 U5499 ( .A(net217232), .ZN(net219494) );
  NAND3_X2 U5500 ( .A1(net217086), .A2(net219494), .A3(net217084), .ZN(
        net216653) );
  INV_X4 U5501 ( .A(net217085), .ZN(net217232) );
  OAI211_X2 U5502 ( .C1(net217232), .C2(net217233), .A(net217231), .B(
        net219976), .ZN(net217228) );
  OAI21_X4 U5503 ( .B1(net215793), .B2(n3650), .A(n3603), .ZN(net215668) );
  XNOR2_X2 U5504 ( .A(n3651), .B(n3603), .ZN(net220293) );
  INV_X4 U5505 ( .A(net215797), .ZN(n3650) );
  INV_X8 U5506 ( .A(net216092), .ZN(net215793) );
  OAI21_X4 U5507 ( .B1(net215793), .B2(net216193), .A(net216192), .ZN(
        net216001) );
  NAND2_X4 U5508 ( .A1(net219781), .A2(net216208), .ZN(net216018) );
  INV_X4 U5509 ( .A(net216018), .ZN(net216207) );
  NAND3_X4 U5510 ( .A1(net216018), .A2(net216019), .A3(net216020), .ZN(
        net215807) );
  OAI21_X4 U5511 ( .B1(net216582), .B2(net216583), .A(net216572), .ZN(
        net219781) );
  NAND3_X2 U5512 ( .A1(net216565), .A2(net216209), .A3(net216566), .ZN(
        net216202) );
  NAND2_X2 U5513 ( .A1(n3652), .A2(n3653), .ZN(net216208) );
  NAND2_X4 U5514 ( .A1(net219781), .A2(net216208), .ZN(net216388) );
  XNOR2_X1 U5515 ( .A(n3654), .B(net216392), .ZN(n3653) );
  INV_X4 U5516 ( .A(net216394), .ZN(n3652) );
  OAI21_X2 U5517 ( .B1(net216582), .B2(net216583), .A(net216572), .ZN(
        net216209) );
  NAND2_X2 U5518 ( .A1(net216584), .A2(net216392), .ZN(net219238) );
  INV_X1 U5519 ( .A(net216392), .ZN(net219237) );
  XNOR2_X2 U5520 ( .A(n3654), .B(net216394), .ZN(net216584) );
  NAND2_X2 U5521 ( .A1(net217631), .A2(net216394), .ZN(net217439) );
  NAND2_X4 U5522 ( .A1(net218061), .A2(net218060), .ZN(net217231) );
  NAND2_X4 U5523 ( .A1(net217085), .A2(net217231), .ZN(net218054) );
  NAND3_X2 U5524 ( .A1(net217231), .A2(net217230), .A3(net217229), .ZN(
        net217086) );
  INV_X4 U5525 ( .A(net218063), .ZN(net218060) );
  INV_X4 U5526 ( .A(n3196), .ZN(net218061) );
  NAND2_X2 U5527 ( .A1(b[5]), .A2(net219055), .ZN(net218063) );
  NAND2_X2 U5528 ( .A1(net218063), .A2(net223531), .ZN(net217085) );
  XNOR2_X2 U5529 ( .A(n3655), .B(net218065), .ZN(net223531) );
  AOI21_X4 U5530 ( .B1(n3656), .B2(n3420), .A(n3657), .ZN(n3655) );
  INV_X8 U5531 ( .A(n3288), .ZN(net218109) );
  NAND2_X4 U5532 ( .A1(n3658), .A2(net220019), .ZN(n3656) );
  NAND2_X2 U5533 ( .A1(net218140), .A2(net217237), .ZN(net218135) );
  OAI21_X4 U5534 ( .B1(net217237), .B2(net217238), .A(n3288), .ZN(net216947)
         );
  NAND3_X1 U5535 ( .A1(net218143), .A2(net218116), .A3(net218115), .ZN(n3658)
         );
  NAND2_X2 U5536 ( .A1(b[9]), .A2(a[11]), .ZN(net215351) );
  INV_X4 U5537 ( .A(net214960), .ZN(net214959) );
  INV_X2 U5538 ( .A(net214961), .ZN(net214954) );
  NAND2_X4 U5539 ( .A1(net212652), .A2(net212649), .ZN(net213006) );
  OAI21_X4 U5540 ( .B1(net213887), .B2(net213888), .A(net213889), .ZN(
        net213588) );
  XNOR2_X2 U5541 ( .A(net213719), .B(net213588), .ZN(net213716) );
  INV_X2 U5542 ( .A(net213588), .ZN(net213586) );
  NOR2_X2 U5543 ( .A1(net213891), .A2(net219539), .ZN(net213888) );
  INV_X4 U5544 ( .A(net213892), .ZN(net213887) );
  NAND2_X2 U5545 ( .A1(n3659), .A2(net213984), .ZN(net213889) );
  NAND2_X4 U5546 ( .A1(net213889), .A2(net213892), .ZN(net213981) );
  INV_X4 U5547 ( .A(net213983), .ZN(n3659) );
  INV_X2 U5548 ( .A(net213891), .ZN(net214172) );
  INV_X4 U5549 ( .A(net220149), .ZN(net214174) );
  NOR2_X4 U5550 ( .A1(net219540), .A2(n3661), .ZN(net219539) );
  NOR2_X4 U5551 ( .A1(net219539), .A2(n3601), .ZN(net214288) );
  INV_X4 U5552 ( .A(n3662), .ZN(n3661) );
  XNOR2_X2 U5553 ( .A(net213989), .B(n3663), .ZN(n3662) );
  NAND2_X4 U5554 ( .A1(net213990), .A2(net213988), .ZN(n3663) );
  NAND2_X4 U5555 ( .A1(net213982), .A2(net213983), .ZN(net213892) );
  INV_X4 U5556 ( .A(net213984), .ZN(net213982) );
  NAND2_X2 U5557 ( .A1(net213989), .A2(net213990), .ZN(n3660) );
  NAND2_X2 U5558 ( .A1(n3660), .A2(net213988), .ZN(net213726) );
  OAI21_X4 U5559 ( .B1(n3664), .B2(net214963), .A(net215332), .ZN(net215217)
         );
  INV_X4 U5560 ( .A(net215217), .ZN(net215216) );
  NOR2_X4 U5561 ( .A1(net214963), .A2(net214964), .ZN(net215114) );
  NAND2_X2 U5562 ( .A1(b[11]), .A2(a[9]), .ZN(net215332) );
  INV_X4 U5563 ( .A(net215332), .ZN(net215329) );
  NAND2_X4 U5564 ( .A1(net215337), .A2(net215338), .ZN(net215331) );
  CLKBUF_X3 U5565 ( .A(net215335), .Z(n3667) );
  NAND3_X4 U5566 ( .A1(net215336), .A2(n3667), .A3(n3666), .ZN(net215330) );
  NAND3_X2 U5567 ( .A1(net215329), .A2(net223718), .A3(net215330), .ZN(
        net214969) );
  INV_X2 U5568 ( .A(n3665), .ZN(n3666) );
  INV_X2 U5569 ( .A(net215337), .ZN(net215336) );
  NAND2_X2 U5570 ( .A1(net219220), .A2(net216094), .ZN(net215797) );
  XNOR2_X1 U5571 ( .A(net216210), .B(net216205), .ZN(net216094) );
  NAND3_X4 U5572 ( .A1(net218271), .A2(net218270), .A3(net218269), .ZN(
        net218216) );
  INV_X8 U5573 ( .A(net220033), .ZN(net218276) );
  NAND2_X4 U5574 ( .A1(net218216), .A2(net218217), .ZN(net218239) );
  NAND2_X4 U5575 ( .A1(net218216), .A2(net218217), .ZN(net218099) );
  NAND2_X4 U5576 ( .A1(net218273), .A2(net218272), .ZN(net218271) );
  NAND2_X2 U5577 ( .A1(net219116), .A2(net217081), .ZN(net216652) );
  INV_X4 U5578 ( .A(net216652), .ZN(net216650) );
  XOR2_X2 U5579 ( .A(net217235), .B(net217082), .Z(net219976) );
  NAND2_X2 U5580 ( .A1(net216941), .A2(net216945), .ZN(net217094) );
  NAND2_X4 U5581 ( .A1(net216941), .A2(net216945), .ZN(net216819) );
  NAND2_X4 U5582 ( .A1(net217230), .A2(net217229), .ZN(net217295) );
  OAI21_X4 U5583 ( .B1(net213586), .B2(n3668), .A(n3673), .ZN(net213233) );
  INV_X2 U5584 ( .A(n3672), .ZN(n3673) );
  INV_X2 U5585 ( .A(net213587), .ZN(n3672) );
  INV_X2 U5586 ( .A(net213589), .ZN(n3668) );
  NAND2_X4 U5587 ( .A1(net213589), .A2(net213587), .ZN(net213719) );
  XNOR2_X2 U5588 ( .A(net213724), .B(net213725), .ZN(n3674) );
  XNOR2_X2 U5589 ( .A(net213724), .B(net213725), .ZN(n3670) );
  INV_X4 U5590 ( .A(net213722), .ZN(n3669) );
  NAND2_X4 U5591 ( .A1(n3671), .A2(net213722), .ZN(net213589) );
  NAND2_X4 U5592 ( .A1(b[1]), .A2(a[1]), .ZN(net217863) );
  OAI21_X1 U5593 ( .B1(net218556), .B2(a[1]), .A(net217863), .ZN(net217433) );
  INV_X4 U5594 ( .A(net217863), .ZN(net218354) );
  NAND2_X4 U5595 ( .A1(net216773), .A2(net216774), .ZN(n3675) );
  NAND2_X4 U5596 ( .A1(net216585), .A2(n3675), .ZN(net216392) );
  NAND2_X4 U5597 ( .A1(net216585), .A2(n3675), .ZN(net216222) );
  INV_X4 U5598 ( .A(net216775), .ZN(net216774) );
  INV_X4 U5599 ( .A(net216776), .ZN(net216773) );
  NAND2_X2 U5600 ( .A1(net216776), .A2(net216775), .ZN(net216226) );
  NAND2_X2 U5601 ( .A1(b[6]), .A2(a[7]), .ZN(net216776) );
  XNOR2_X2 U5602 ( .A(net215339), .B(net214877), .ZN(net215337) );
  NAND2_X2 U5603 ( .A1(net217550), .A2(net215210), .ZN(net217299) );
  NOR2_X4 U5604 ( .A1(net215209), .A2(net215210), .ZN(net214964) );
  AOI21_X4 U5605 ( .B1(n3683), .B2(n3685), .A(net215216), .ZN(net214967) );
  INV_X2 U5606 ( .A(n3684), .ZN(n3685) );
  INV_X4 U5607 ( .A(net215215), .ZN(n3684) );
  INV_X4 U5608 ( .A(net215446), .ZN(n3677) );
  OAI21_X2 U5609 ( .B1(n3677), .B2(n3676), .A(net215445), .ZN(net215214) );
  INV_X4 U5610 ( .A(net215447), .ZN(n3676) );
  NAND2_X4 U5611 ( .A1(net215215), .A2(net215445), .ZN(net215566) );
  INV_X4 U5612 ( .A(net215568), .ZN(n3679) );
  NAND2_X4 U5613 ( .A1(n3678), .A2(net215568), .ZN(net215445) );
  INV_X4 U5614 ( .A(n3427), .ZN(n3678) );
  OAI21_X4 U5615 ( .B1(n3680), .B2(n3681), .A(net215672), .ZN(net215446) );
  NAND2_X2 U5616 ( .A1(net215446), .A2(net215447), .ZN(net215565) );
  INV_X4 U5617 ( .A(net215673), .ZN(n3681) );
  INV_X1 U5618 ( .A(net215674), .ZN(n3680) );
  NAND2_X4 U5619 ( .A1(net215672), .A2(net215447), .ZN(net215770) );
  INV_X4 U5620 ( .A(net215773), .ZN(n3682) );
  XNOR2_X2 U5621 ( .A(net215775), .B(net215776), .ZN(n3686) );
  AOI21_X2 U5622 ( .B1(net214831), .B2(net214832), .A(net215081), .ZN(n3687)
         );
  INV_X4 U5623 ( .A(net215081), .ZN(net220181) );
  INV_X4 U5624 ( .A(net215082), .ZN(net215078) );
  NAND2_X2 U5625 ( .A1(b[16]), .A2(a[5]), .ZN(net215076) );
  NAND2_X2 U5626 ( .A1(net214831), .A2(net214832), .ZN(net214571) );
  XNOR2_X2 U5627 ( .A(n3688), .B(net214831), .ZN(net215300) );
  AOI21_X4 U5628 ( .B1(net212642), .B2(net219746), .A(net212644), .ZN(
        net212640) );
  NOR3_X4 U5629 ( .A1(n3689), .A2(n3692), .A3(n3690), .ZN(net216582) );
  INV_X4 U5630 ( .A(net216660), .ZN(n3690) );
  INV_X4 U5631 ( .A(net216577), .ZN(n3695) );
  INV_X2 U5632 ( .A(net216578), .ZN(n3694) );
  INV_X2 U5633 ( .A(n3694), .ZN(net219847) );
  INV_X2 U5634 ( .A(net216579), .ZN(net216658) );
  INV_X4 U5635 ( .A(net216761), .ZN(net216657) );
  NAND2_X2 U5636 ( .A1(net216657), .A2(net219526), .ZN(net216576) );
  INV_X4 U5637 ( .A(net219526), .ZN(net216762) );
  NAND2_X4 U5638 ( .A1(net216762), .A2(net216761), .ZN(n3693) );
  NAND2_X4 U5639 ( .A1(n3696), .A2(net219238), .ZN(net216572) );
  INV_X4 U5640 ( .A(net216584), .ZN(net219236) );
  NAND2_X4 U5641 ( .A1(net216836), .A2(net216660), .ZN(net216759) );
  NAND2_X4 U5642 ( .A1(n3697), .A2(net217088), .ZN(net216651) );
  OAI21_X4 U5643 ( .B1(net216649), .B2(net216650), .A(net216651), .ZN(
        net216647) );
  XNOR2_X1 U5644 ( .A(net217092), .B(net217091), .ZN(n3697) );
  NAND2_X4 U5645 ( .A1(net216935), .A2(net216934), .ZN(net219641) );
  NAND2_X4 U5646 ( .A1(net215061), .A2(n3701), .ZN(net214545) );
  INV_X4 U5647 ( .A(net215062), .ZN(n3701) );
  NAND2_X4 U5648 ( .A1(n3698), .A2(net214786), .ZN(net214546) );
  OAI21_X4 U5649 ( .B1(n3699), .B2(n3700), .A(net214983), .ZN(n3698) );
  INV_X4 U5650 ( .A(net215058), .ZN(n3699) );
  OAI21_X2 U5651 ( .B1(n3699), .B2(n3700), .A(net214983), .ZN(net214785) );
  NAND2_X4 U5652 ( .A1(n3702), .A2(net215062), .ZN(net214786) );
  XNOR2_X2 U5653 ( .A(net215058), .B(n3703), .ZN(net215275) );
  NAND2_X2 U5654 ( .A1(net213406), .A2(net213407), .ZN(net213237) );
  INV_X4 U5655 ( .A(net213405), .ZN(net213407) );
  INV_X4 U5656 ( .A(net213406), .ZN(net213404) );
  NAND2_X2 U5657 ( .A1(a[8]), .A2(b[19]), .ZN(net213405) );
  NAND2_X4 U5658 ( .A1(net213404), .A2(net213405), .ZN(net213239) );
  NAND2_X2 U5659 ( .A1(a[7]), .A2(b[20]), .ZN(net213400) );
  NAND3_X2 U5660 ( .A1(n3707), .A2(net218135), .A3(net218136), .ZN(net217229)
         );
  INV_X4 U5661 ( .A(net218137), .ZN(n3707) );
  OAI211_X4 U5662 ( .C1(n3704), .C2(n3705), .A(net218042), .B(net218057), .ZN(
        net217230) );
  NAND2_X2 U5663 ( .A1(net218058), .A2(net218059), .ZN(n3705) );
  INV_X4 U5664 ( .A(net218043), .ZN(n3704) );
  NOR2_X4 U5665 ( .A1(n3704), .A2(n3706), .ZN(net218124) );
  OAI21_X4 U5666 ( .B1(n3708), .B2(net218139), .A(net218137), .ZN(net218057)
         );
  INV_X4 U5667 ( .A(net218042), .ZN(n3706) );
  NAND2_X4 U5668 ( .A1(net218058), .A2(net218059), .ZN(net218041) );
  OAI21_X4 U5669 ( .B1(n3706), .B2(net218178), .A(net218043), .ZN(net218132)
         );
  NAND2_X4 U5670 ( .A1(net216844), .A2(net216929), .ZN(net216660) );
  OAI21_X4 U5671 ( .B1(n3709), .B2(n3710), .A(net216839), .ZN(net216577) );
  NAND3_X1 U5672 ( .A1(net216577), .A2(net219847), .A3(net216579), .ZN(
        net216574) );
  NAND3_X2 U5673 ( .A1(net216579), .A2(net219847), .A3(net216577), .ZN(
        net216836) );
  INV_X4 U5674 ( .A(net216840), .ZN(n3710) );
  INV_X1 U5675 ( .A(n3299), .ZN(n3709) );
  NAND2_X2 U5676 ( .A1(n3711), .A2(net217070), .ZN(net216578) );
  INV_X4 U5677 ( .A(net217071), .ZN(n3711) );
  NAND2_X2 U5678 ( .A1(n3711), .A2(net216987), .ZN(net216985) );
  INV_X1 U5679 ( .A(net216844), .ZN(net216843) );
  INV_X4 U5680 ( .A(net216929), .ZN(net216842) );
  NAND2_X4 U5681 ( .A1(net214720), .A2(net214721), .ZN(net214817) );
  NAND2_X4 U5682 ( .A1(net215324), .A2(n3712), .ZN(net214856) );
  INV_X4 U5683 ( .A(net215325), .ZN(n3712) );
  INV_X4 U5684 ( .A(net215324), .ZN(n3713) );
  NAND2_X4 U5685 ( .A1(n3713), .A2(net215325), .ZN(net215219) );
  XNOR2_X2 U5686 ( .A(net215218), .B(net215322), .ZN(net215318) );
  NAND2_X4 U5687 ( .A1(n3714), .A2(n3327), .ZN(net214727) );
  XNOR2_X2 U5688 ( .A(net215072), .B(net215073), .ZN(n3714) );
  NAND2_X4 U5689 ( .A1(net215295), .A2(net215296), .ZN(net214804) );
  NAND2_X4 U5690 ( .A1(net214804), .A2(net214730), .ZN(net215287) );
  OAI21_X4 U5691 ( .B1(net219358), .B2(net217285), .A(n3715), .ZN(net217109)
         );
  NAND4_X2 U5692 ( .A1(net217291), .A2(net217293), .A3(net217292), .A4(
        net217294), .ZN(net218101) );
  NAND2_X4 U5693 ( .A1(net218105), .A2(net218106), .ZN(net217290) );
  INV_X1 U5694 ( .A(net219358), .ZN(net217283) );
  NAND2_X4 U5695 ( .A1(net217284), .A2(net217285), .ZN(n3715) );
  INV_X4 U5696 ( .A(net217285), .ZN(net217282) );
  NAND3_X2 U5697 ( .A1(net217106), .A2(net219368), .A3(n3715), .ZN(net217281)
         );
  NAND2_X2 U5698 ( .A1(net217294), .A2(net217293), .ZN(net217287) );
  NAND2_X4 U5699 ( .A1(n3716), .A2(net214834), .ZN(net214831) );
  NAND2_X4 U5700 ( .A1(n3718), .A2(net215468), .ZN(n3716) );
  OAI21_X4 U5701 ( .B1(n3719), .B2(n3720), .A(n3724), .ZN(n3718) );
  INV_X4 U5702 ( .A(n3723), .ZN(n3724) );
  INV_X4 U5703 ( .A(net215471), .ZN(n3723) );
  AOI21_X2 U5704 ( .B1(net215675), .B2(net215478), .A(n3723), .ZN(net215530)
         );
  OAI21_X4 U5705 ( .B1(n3721), .B2(net220410), .A(n3722), .ZN(n3720) );
  NAND3_X4 U5706 ( .A1(net215475), .A2(n3725), .A3(net215477), .ZN(n3722) );
  CLKBUF_X3 U5707 ( .A(net215476), .Z(n3725) );
  INV_X4 U5708 ( .A(net215478), .ZN(n3719) );
  NAND2_X4 U5709 ( .A1(net215308), .A2(net215307), .ZN(net214832) );
  INV_X4 U5710 ( .A(net223908), .ZN(net215308) );
  NAND2_X4 U5711 ( .A1(net223908), .A2(n3717), .ZN(net214569) );
  INV_X4 U5712 ( .A(net215307), .ZN(n3717) );
  NAND2_X4 U5713 ( .A1(n3727), .A2(n3726), .ZN(net217262) );
  INV_X4 U5714 ( .A(net218157), .ZN(n3726) );
  NAND2_X4 U5715 ( .A1(n3727), .A2(n3726), .ZN(net220022) );
  INV_X4 U5716 ( .A(net218156), .ZN(n3727) );
  NAND3_X4 U5717 ( .A1(net218219), .A2(net218220), .A3(net218221), .ZN(
        net218098) );
  INV_X4 U5718 ( .A(net218174), .ZN(net218221) );
  NAND2_X4 U5719 ( .A1(net218173), .A2(net218174), .ZN(net218094) );
  NAND2_X2 U5720 ( .A1(net218550), .A2(a[5]), .ZN(net218174) );
  NAND2_X4 U5721 ( .A1(n3730), .A2(net215357), .ZN(net214960) );
  INV_X4 U5722 ( .A(n3733), .ZN(n3730) );
  XNOR2_X2 U5723 ( .A(n3731), .B(net215360), .ZN(n3733) );
  INV_X4 U5724 ( .A(net215357), .ZN(n3728) );
  NAND2_X2 U5725 ( .A1(n3735), .A2(net215112), .ZN(net214864) );
  INV_X4 U5726 ( .A(net215111), .ZN(n3735) );
  NAND2_X4 U5727 ( .A1(n3734), .A2(net215111), .ZN(net214968) );
  INV_X4 U5728 ( .A(net215112), .ZN(n3734) );
  XNOR2_X2 U5729 ( .A(net216763), .B(n3740), .ZN(net219526) );
  INV_X4 U5730 ( .A(n3743), .ZN(n3741) );
  INV_X4 U5731 ( .A(n3744), .ZN(n3739) );
  NAND3_X2 U5732 ( .A1(n3746), .A2(n3739), .A3(net219497), .ZN(net216927) );
  NAND3_X2 U5733 ( .A1(n3738), .A2(net219497), .A3(n3746), .ZN(n3737) );
  INV_X4 U5734 ( .A(net216979), .ZN(n3742) );
  XNOR2_X2 U5735 ( .A(net216978), .B(n3742), .ZN(n3745) );
  NAND2_X2 U5736 ( .A1(n3746), .A2(net216587), .ZN(n3743) );
  NAND2_X1 U5737 ( .A1(n3743), .A2(n3744), .ZN(net216928) );
  XNOR2_X2 U5738 ( .A(n3745), .B(net216835), .ZN(n3744) );
  NAND3_X2 U5739 ( .A1(n3736), .A2(net216226), .A3(n3737), .ZN(net216585) );
  OAI21_X4 U5740 ( .B1(n3748), .B2(n3747), .A(n3751), .ZN(net213238) );
  INV_X2 U5741 ( .A(n3750), .ZN(n3751) );
  INV_X2 U5742 ( .A(net213592), .ZN(n3750) );
  INV_X2 U5743 ( .A(net213594), .ZN(n3747) );
  NAND2_X4 U5744 ( .A1(net213594), .A2(net213592), .ZN(n3749) );
  XNOR2_X2 U5745 ( .A(net213593), .B(n3749), .ZN(net213711) );
  NAND2_X4 U5746 ( .A1(net212740), .A2(net212739), .ZN(net212641) );
  OAI21_X4 U5747 ( .B1(n3308), .B2(n3752), .A(net216283), .ZN(net216282) );
  XNOR2_X1 U5748 ( .A(net216783), .B(net216782), .ZN(n3752) );
  NAND2_X2 U5749 ( .A1(n3753), .A2(net213411), .ZN(net213232) );
  INV_X4 U5750 ( .A(net213410), .ZN(n3753) );
  NAND2_X4 U5751 ( .A1(net213409), .A2(net213410), .ZN(net213234) );
  INV_X4 U5752 ( .A(net213411), .ZN(net213409) );
  NAND2_X4 U5753 ( .A1(n3754), .A2(net218281), .ZN(net218100) );
  NAND2_X4 U5754 ( .A1(net218097), .A2(net218100), .ZN(net218238) );
  XNOR2_X2 U5755 ( .A(net218284), .B(net218285), .ZN(n3754) );
  OAI21_X4 U5756 ( .B1(n3755), .B2(n3756), .A(net215342), .ZN(net214877) );
  INV_X2 U5757 ( .A(net214877), .ZN(net215211) );
  AOI21_X2 U5758 ( .B1(net215344), .B2(net219978), .A(n3757), .ZN(n3756) );
  INV_X4 U5759 ( .A(net215346), .ZN(n3757) );
  NAND2_X4 U5760 ( .A1(net219978), .A2(net215344), .ZN(net215583) );
  INV_X4 U5761 ( .A(net215343), .ZN(net215784) );
  NAND3_X2 U5762 ( .A1(net215782), .A2(net215783), .A3(net215784), .ZN(
        net215777) );
  XNOR2_X2 U5763 ( .A(net215586), .B(net215792), .ZN(net215343) );
  NAND2_X2 U5764 ( .A1(net223270), .A2(net223271), .ZN(net215792) );
  INV_X4 U5765 ( .A(net215347), .ZN(n3755) );
  INV_X4 U5766 ( .A(net214846), .ZN(net223412) );
  NOR2_X4 U5767 ( .A1(n3759), .A2(n6349), .ZN(n3758) );
  INV_X4 U5768 ( .A(n3758), .ZN(n6532) );
  AND2_X2 U5769 ( .A1(a[19]), .A2(b[4]), .ZN(n3759) );
  OAI21_X2 U5770 ( .B1(n5926), .B2(n6036), .A(n6035), .ZN(n6172) );
  INV_X2 U5771 ( .A(n4410), .ZN(n4411) );
  OAI21_X2 U5772 ( .B1(n7261), .B2(net212881), .A(n7260), .ZN(n7408) );
  INV_X2 U5773 ( .A(n5288), .ZN(n5291) );
  NAND2_X4 U5774 ( .A1(n4714), .A2(net220022), .ZN(net217258) );
  NAND2_X4 U5775 ( .A1(net217261), .A2(net220022), .ZN(net217260) );
  AND2_X2 U5776 ( .A1(n7140), .A2(n7139), .ZN(n3760) );
  NAND2_X4 U5777 ( .A1(a[23]), .A2(b[5]), .ZN(n7140) );
  INV_X2 U5778 ( .A(n4121), .ZN(n4016) );
  NAND2_X4 U5779 ( .A1(n5107), .A2(n5106), .ZN(n5246) );
  NAND2_X4 U5780 ( .A1(n6233), .A2(n3871), .ZN(n6397) );
  XNOR2_X2 U5781 ( .A(n6740), .B(n6553), .ZN(n3761) );
  INV_X4 U5782 ( .A(n3761), .ZN(n6555) );
  NAND2_X2 U5783 ( .A1(net218238), .A2(n3863), .ZN(n3809) );
  INV_X2 U5784 ( .A(net218244), .ZN(net218263) );
  BUF_X4 U5785 ( .A(net218115), .Z(net224032) );
  OAI21_X2 U5786 ( .B1(net218260), .B2(net218261), .A(net218240), .ZN(n3839)
         );
  XNOR2_X2 U5787 ( .A(n5563), .B(n5561), .ZN(n3762) );
  NAND2_X4 U5788 ( .A1(n5898), .A2(n5620), .ZN(n5561) );
  NAND2_X4 U5789 ( .A1(n3764), .A2(n5915), .ZN(net215776) );
  NAND2_X1 U5790 ( .A1(n4029), .A2(n4007), .ZN(n3763) );
  INV_X4 U5791 ( .A(n5957), .ZN(n5811) );
  INV_X2 U5792 ( .A(net212470), .ZN(net212468) );
  NAND2_X4 U5793 ( .A1(n5971), .A2(net215294), .ZN(net224078) );
  INV_X1 U5794 ( .A(n3882), .ZN(n3807) );
  XNOR2_X2 U5795 ( .A(n6614), .B(n6613), .ZN(n3765) );
  OAI22_X4 U5796 ( .A1(n5770), .A2(n5769), .B1(net220410), .B2(n5715), .ZN(
        n5585) );
  INV_X2 U5797 ( .A(net213553), .ZN(net214024) );
  OAI21_X1 U5798 ( .B1(n3219), .B2(net213766), .A(net213553), .ZN(net213763)
         );
  INV_X4 U5799 ( .A(net212653), .ZN(net219657) );
  NAND2_X2 U5800 ( .A1(n7292), .A2(n7291), .ZN(n3767) );
  NAND2_X4 U5801 ( .A1(n7140), .A2(n7139), .ZN(n7291) );
  NAND2_X4 U5802 ( .A1(n7234), .A2(n7233), .ZN(n7235) );
  XNOR2_X2 U5803 ( .A(net213005), .B(net213006), .ZN(n3768) );
  NAND2_X4 U5804 ( .A1(n3781), .A2(n7194), .ZN(net212649) );
  XNOR2_X2 U5805 ( .A(net214610), .B(net214611), .ZN(n3769) );
  NAND2_X4 U5806 ( .A1(n3845), .A2(n3853), .ZN(net214611) );
  OAI21_X4 U5807 ( .B1(n4970), .B2(n4969), .A(n4968), .ZN(n3770) );
  NAND2_X4 U5808 ( .A1(n4927), .A2(n3794), .ZN(n4968) );
  XNOR2_X2 U5809 ( .A(n6801), .B(n6802), .ZN(n3771) );
  NAND2_X4 U5810 ( .A1(n6692), .A2(n3918), .ZN(net213576) );
  NAND2_X2 U5811 ( .A1(n7172), .A2(n7171), .ZN(n7500) );
  INV_X2 U5812 ( .A(n6223), .ZN(n6224) );
  NAND2_X4 U5813 ( .A1(n7340), .A2(n7339), .ZN(n7513) );
  XNOR2_X2 U5814 ( .A(net212881), .B(n7152), .ZN(n3772) );
  INV_X4 U5815 ( .A(n3772), .ZN(n7154) );
  NAND2_X4 U5816 ( .A1(n5341), .A2(n5630), .ZN(n5297) );
  INV_X8 U5817 ( .A(n6028), .ZN(n5959) );
  NAND2_X4 U5818 ( .A1(n3376), .A2(n6611), .ZN(n6667) );
  XNOR2_X2 U5819 ( .A(n6610), .B(n3937), .ZN(n6611) );
  OAI21_X4 U5820 ( .B1(net214711), .B2(net214710), .A(n6301), .ZN(n6494) );
  XOR2_X2 U5821 ( .A(net215581), .B(net215582), .Z(n3773) );
  NAND2_X4 U5822 ( .A1(net215347), .A2(net215342), .ZN(net215581) );
  NAND2_X4 U5823 ( .A1(net215583), .A2(net215346), .ZN(net215582) );
  XOR2_X2 U5824 ( .A(net218054), .B(net217295), .Z(n3774) );
  INV_X2 U5825 ( .A(n5373), .ZN(n5376) );
  XNOR2_X2 U5826 ( .A(n3776), .B(n4801), .ZN(n3775) );
  INV_X4 U5827 ( .A(n3775), .ZN(n4803) );
  INV_X2 U5828 ( .A(n5888), .ZN(n3777) );
  NAND2_X4 U5829 ( .A1(n4994), .A2(net216794), .ZN(n5099) );
  INV_X2 U5830 ( .A(net216794), .ZN(net216795) );
  AOI21_X2 U5831 ( .B1(n3416), .B2(n5211), .A(n5210), .ZN(n3778) );
  NAND2_X2 U5832 ( .A1(n5208), .A2(n5207), .ZN(n5211) );
  XNOR2_X2 U5833 ( .A(net212906), .B(n7246), .ZN(n3779) );
  INV_X8 U5834 ( .A(n4082), .ZN(n4380) );
  INV_X2 U5835 ( .A(n5571), .ZN(n5572) );
  NAND2_X1 U5836 ( .A1(n5435), .A2(n5571), .ZN(n5307) );
  OAI21_X2 U5837 ( .B1(n5436), .B2(n5568), .A(n5571), .ZN(n5437) );
  AOI21_X2 U5838 ( .B1(n5570), .B2(n5569), .A(n5568), .ZN(n5573) );
  OAI21_X4 U5839 ( .B1(n5648), .B2(n5647), .A(n5646), .ZN(n3780) );
  NAND2_X4 U5840 ( .A1(n4983), .A2(n5092), .ZN(n4903) );
  XNOR2_X2 U5841 ( .A(n3476), .B(net213012), .ZN(n3781) );
  OAI21_X4 U5842 ( .B1(net217288), .B2(net217287), .A(net219864), .ZN(n3782)
         );
  XNOR2_X2 U5843 ( .A(n6368), .B(n6367), .ZN(n3783) );
  OAI21_X2 U5844 ( .B1(n7493), .B2(n7492), .A(n7491), .ZN(n7496) );
  INV_X2 U5845 ( .A(n7171), .ZN(n7169) );
  XNOR2_X2 U5846 ( .A(n5850), .B(n5849), .ZN(n3784) );
  AOI21_X2 U5847 ( .B1(n5848), .B2(n5895), .A(n5847), .ZN(n5849) );
  XNOR2_X1 U5848 ( .A(n3858), .B(net216096), .ZN(n3785) );
  INV_X8 U5849 ( .A(n5416), .ZN(n5419) );
  OAI21_X2 U5850 ( .B1(n3307), .B2(n3962), .A(n5803), .ZN(n3786) );
  AND3_X4 U5851 ( .A1(net215777), .A2(net215583), .A3(n5690), .ZN(n3787) );
  INV_X4 U5852 ( .A(n3787), .ZN(n5915) );
  NAND2_X4 U5853 ( .A1(n7484), .A2(n7482), .ZN(n7313) );
  NAND2_X4 U5854 ( .A1(n7312), .A2(n7311), .ZN(n7482) );
  NAND2_X4 U5855 ( .A1(n4052), .A2(net218282), .ZN(net223819) );
  INV_X8 U5856 ( .A(net212902), .ZN(net212906) );
  NAND2_X4 U5857 ( .A1(net215320), .A2(n5963), .ZN(net215224) );
  CLKBUF_X2 U5858 ( .A(n5935), .Z(n3788) );
  NAND2_X2 U5859 ( .A1(n6681), .A2(n6685), .ZN(n6435) );
  NAND2_X4 U5860 ( .A1(net213577), .A2(net213736), .ZN(net213997) );
  NAND2_X4 U5861 ( .A1(n6688), .A2(n6687), .ZN(n6690) );
  INV_X2 U5862 ( .A(net214385), .ZN(net214387) );
  NAND2_X1 U5863 ( .A1(n6334), .A2(n6335), .ZN(n6182) );
  NAND2_X4 U5864 ( .A1(n3860), .A2(n3861), .ZN(n3858) );
  NAND2_X2 U5865 ( .A1(net216095), .A2(net216097), .ZN(n3860) );
  NAND2_X4 U5866 ( .A1(n7761), .A2(n7760), .ZN(n7524) );
  NAND2_X4 U5867 ( .A1(net212646), .A2(net219679), .ZN(net212134) );
  XNOR2_X2 U5868 ( .A(n7590), .B(n7591), .ZN(n3789) );
  INV_X4 U5869 ( .A(n3789), .ZN(n7522) );
  NAND2_X1 U5870 ( .A1(a[15]), .A2(b[15]), .ZN(n7589) );
  INV_X2 U5871 ( .A(n7589), .ZN(n7591) );
  NAND3_X2 U5872 ( .A1(net211934), .A2(net211935), .A3(n3355), .ZN(result[31])
         );
  OAI21_X4 U5873 ( .B1(net212099), .B2(net218614), .A(net212102), .ZN(
        net211935) );
  AND2_X2 U5874 ( .A1(net220298), .A2(net212394), .ZN(n3821) );
  INV_X4 U5875 ( .A(net211935), .ZN(net211942) );
  INV_X1 U5876 ( .A(net223617), .ZN(net223581) );
  NAND3_X2 U5877 ( .A1(net212685), .A2(net212686), .A3(net212687), .ZN(
        net212404) );
  NAND2_X4 U5878 ( .A1(net223484), .A2(net212691), .ZN(net212685) );
  XNOR2_X2 U5879 ( .A(net214840), .B(n6239), .ZN(n3790) );
  CLKBUF_X2 U5880 ( .A(n5077), .Z(n3791) );
  NAND2_X4 U5881 ( .A1(n3202), .A2(n4917), .ZN(n5077) );
  NAND2_X1 U5882 ( .A1(n6089), .A2(n6428), .ZN(n5985) );
  XNOR2_X2 U5883 ( .A(n6584), .B(n6585), .ZN(n3792) );
  XNOR2_X2 U5884 ( .A(n5278), .B(n5277), .ZN(n3793) );
  XNOR2_X2 U5885 ( .A(n4923), .B(n4922), .ZN(n3794) );
  NAND2_X4 U5886 ( .A1(n4840), .A2(n5074), .ZN(n4922) );
  XNOR2_X2 U5887 ( .A(n5266), .B(net216388), .ZN(n3795) );
  NAND2_X4 U5888 ( .A1(n5141), .A2(n5292), .ZN(n5142) );
  NAND2_X4 U5889 ( .A1(n5295), .A2(n5538), .ZN(n5143) );
  NAND3_X2 U5890 ( .A1(a[0]), .A2(b[11]), .A3(n4934), .ZN(n5288) );
  NAND2_X2 U5891 ( .A1(n6219), .A2(n6220), .ZN(net214434) );
  NAND3_X2 U5892 ( .A1(n7375), .A2(a[0]), .A3(b[28]), .ZN(net212412) );
  XNOR2_X2 U5893 ( .A(n7263), .B(net213111), .ZN(n7144) );
  XNOR2_X2 U5894 ( .A(n5818), .B(net215593), .ZN(n3796) );
  INV_X4 U5895 ( .A(n5130), .ZN(n3813) );
  INV_X4 U5896 ( .A(net216944), .ZN(net217236) );
  XNOR2_X2 U5897 ( .A(n6797), .B(n6798), .ZN(n3797) );
  INV_X2 U5898 ( .A(n5394), .ZN(n5395) );
  INV_X2 U5899 ( .A(n6786), .ZN(n6575) );
  NAND2_X4 U5900 ( .A1(n6314), .A2(n6313), .ZN(n6513) );
  NAND2_X4 U5901 ( .A1(n6773), .A2(n6774), .ZN(net213866) );
  NAND2_X4 U5902 ( .A1(n3798), .A2(n3799), .ZN(n3801) );
  NAND2_X4 U5903 ( .A1(n3800), .A2(n3801), .ZN(n6223) );
  INV_X4 U5904 ( .A(n6221), .ZN(n3798) );
  INV_X2 U5905 ( .A(net214603), .ZN(n3799) );
  INV_X4 U5906 ( .A(net217242), .ZN(net218808) );
  NAND2_X4 U5907 ( .A1(n6080), .A2(n6079), .ZN(n6151) );
  OAI21_X4 U5908 ( .B1(net216206), .B2(net216207), .A(n3862), .ZN(net216205)
         );
  INV_X4 U5909 ( .A(n5617), .ZN(n5562) );
  INV_X4 U5910 ( .A(n5629), .ZN(n5543) );
  NAND2_X4 U5911 ( .A1(net217259), .A2(n4798), .ZN(n4124) );
  OAI21_X4 U5912 ( .B1(n3309), .B2(n5794), .A(n5938), .ZN(n5939) );
  INV_X1 U5913 ( .A(n7553), .ZN(n7555) );
  NAND2_X2 U5914 ( .A1(net214846), .A2(n6234), .ZN(n3803) );
  NAND2_X4 U5915 ( .A1(net223412), .A2(n3802), .ZN(n3804) );
  NAND2_X4 U5916 ( .A1(n3803), .A2(n3804), .ZN(n6236) );
  INV_X4 U5917 ( .A(n6234), .ZN(n3802) );
  NAND2_X4 U5918 ( .A1(net214586), .A2(n6397), .ZN(n6234) );
  INV_X4 U5919 ( .A(n6400), .ZN(n6402) );
  INV_X4 U5920 ( .A(n3769), .ZN(n6379) );
  INV_X2 U5921 ( .A(n5903), .ZN(n5829) );
  NAND2_X2 U5922 ( .A1(n5902), .A2(n3989), .ZN(n5830) );
  INV_X2 U5923 ( .A(n3878), .ZN(n6695) );
  NAND2_X4 U5924 ( .A1(n6232), .A2(n6231), .ZN(net214586) );
  INV_X2 U5925 ( .A(n6680), .ZN(n6487) );
  NOR2_X4 U5926 ( .A1(net218145), .A2(net218147), .ZN(net218233) );
  NAND3_X2 U5927 ( .A1(n5521), .A2(n5523), .A3(n5522), .ZN(n5350) );
  NAND2_X4 U5928 ( .A1(n7332), .A2(n7331), .ZN(n7505) );
  NAND2_X2 U5929 ( .A1(net212792), .A2(n7328), .ZN(n7329) );
  NAND2_X4 U5930 ( .A1(n6601), .A2(n6602), .ZN(n6678) );
  NAND2_X4 U5931 ( .A1(n3769), .A2(n6381), .ZN(n6710) );
  INV_X4 U5932 ( .A(n5485), .ZN(n5378) );
  INV_X1 U5933 ( .A(net214152), .ZN(net214145) );
  NAND2_X4 U5934 ( .A1(n6068), .A2(n6067), .ZN(n6154) );
  INV_X4 U5935 ( .A(n5825), .ZN(n5827) );
  INV_X2 U5936 ( .A(net223586), .ZN(net212114) );
  NAND2_X4 U5937 ( .A1(n6379), .A2(n6380), .ZN(n6712) );
  NAND2_X4 U5938 ( .A1(n5585), .A2(n5584), .ZN(n5764) );
  NAND2_X4 U5939 ( .A1(n5439), .A2(n5440), .ZN(n5581) );
  NAND2_X4 U5940 ( .A1(n5581), .A2(n5579), .ZN(net215475) );
  INV_X4 U5941 ( .A(n5146), .ZN(n5144) );
  NAND3_X2 U5942 ( .A1(n5522), .A2(n5523), .A3(n5521), .ZN(n5524) );
  NAND2_X1 U5943 ( .A1(n3844), .A2(n3845), .ZN(n3847) );
  INV_X4 U5944 ( .A(n3418), .ZN(n6785) );
  NAND2_X1 U5945 ( .A1(n3953), .A2(n6305), .ZN(n3805) );
  CLKBUF_X3 U5946 ( .A(n5355), .Z(n3806) );
  NAND2_X4 U5947 ( .A1(n4899), .A2(n4900), .ZN(n4983) );
  NAND2_X4 U5948 ( .A1(n5347), .A2(n5346), .ZN(n5405) );
  INV_X4 U5949 ( .A(net219641), .ZN(net216645) );
  NAND2_X4 U5950 ( .A1(n5678), .A2(n5679), .ZN(n5773) );
  BUF_X4 U5951 ( .A(n5904), .Z(n3989) );
  INV_X2 U5952 ( .A(n5504), .ZN(n5502) );
  NAND2_X4 U5953 ( .A1(n5886), .A2(n6015), .ZN(n5973) );
  NAND2_X4 U5954 ( .A1(net215478), .A2(net215471), .ZN(n5722) );
  NAND2_X4 U5955 ( .A1(n5123), .A2(net216571), .ZN(net216565) );
  INV_X4 U5956 ( .A(n7338), .ZN(n7340) );
  INV_X2 U5957 ( .A(n7490), .ZN(n7493) );
  OAI21_X1 U5958 ( .B1(n7419), .B2(n7418), .A(n7417), .ZN(n7466) );
  NAND2_X4 U5959 ( .A1(n5655), .A2(n5654), .ZN(n5784) );
  INV_X2 U5960 ( .A(n5493), .ZN(n5370) );
  NAND2_X4 U5961 ( .A1(net214456), .A2(net214457), .ZN(n6490) );
  INV_X4 U5962 ( .A(n7234), .ZN(n3926) );
  INV_X8 U5963 ( .A(n7111), .ZN(n7234) );
  OAI21_X4 U5964 ( .B1(net212927), .B2(net212928), .A(net219674), .ZN(n3882)
         );
  INV_X4 U5965 ( .A(n7542), .ZN(n7544) );
  NAND2_X2 U5966 ( .A1(n6725), .A2(n3203), .ZN(n6566) );
  NAND2_X4 U5967 ( .A1(net214331), .A2(net214332), .ZN(net213556) );
  INV_X2 U5968 ( .A(n5071), .ZN(n3965) );
  NAND2_X1 U5969 ( .A1(n4792), .A2(n4150), .ZN(n4143) );
  NAND2_X4 U5970 ( .A1(n4150), .A2(n4792), .ZN(n4154) );
  INV_X4 U5971 ( .A(n3875), .ZN(n5420) );
  NAND2_X4 U5972 ( .A1(n5153), .A2(n5154), .ZN(n5195) );
  NAND2_X4 U5973 ( .A1(b[9]), .A2(a[9]), .ZN(net215799) );
  OAI21_X2 U5974 ( .B1(net216198), .B2(n5395), .A(net216200), .ZN(n5397) );
  AOI21_X2 U5975 ( .B1(n5913), .B2(n5914), .A(n5912), .ZN(n5916) );
  NAND2_X4 U5976 ( .A1(net218212), .A2(net219965), .ZN(net218106) );
  NAND2_X4 U5977 ( .A1(n5025), .A2(n5024), .ZN(n5212) );
  NAND2_X2 U5978 ( .A1(net213374), .A2(net213373), .ZN(n6970) );
  NAND2_X2 U5979 ( .A1(n5921), .A2(n5920), .ZN(n5788) );
  NAND3_X4 U5980 ( .A1(a[10]), .A2(net216958), .A3(net218548), .ZN(n5104) );
  NAND2_X4 U5981 ( .A1(n5382), .A2(n5381), .ZN(n5643) );
  XNOR2_X1 U5982 ( .A(n4732), .B(n4733), .ZN(n3958) );
  INV_X4 U5983 ( .A(n3946), .ZN(n3808) );
  NAND2_X4 U5984 ( .A1(b[30]), .A2(a[1]), .ZN(n7693) );
  NAND2_X4 U5985 ( .A1(b[14]), .A2(a[1]), .ZN(n5569) );
  NAND2_X4 U5986 ( .A1(b[15]), .A2(a[1]), .ZN(n5440) );
  NAND2_X2 U5987 ( .A1(n4122), .A2(n4121), .ZN(n4103) );
  NAND2_X4 U5988 ( .A1(net216932), .A2(net216587), .ZN(n4819) );
  INV_X2 U5989 ( .A(net217075), .ZN(net217077) );
  NAND2_X4 U5990 ( .A1(n6732), .A2(n6731), .ZN(net213851) );
  INV_X8 U5991 ( .A(net220099), .ZN(net212951) );
  NAND2_X1 U5992 ( .A1(n6767), .A2(n6766), .ZN(n6763) );
  INV_X4 U5993 ( .A(n5351), .ZN(n5353) );
  NAND2_X4 U5994 ( .A1(n5135), .A2(n5136), .ZN(n5538) );
  NAND2_X4 U5995 ( .A1(n6695), .A2(n6885), .ZN(n6584) );
  NAND2_X4 U5996 ( .A1(n3353), .A2(n6583), .ZN(n6885) );
  NAND2_X4 U5997 ( .A1(n5133), .A2(n5134), .ZN(n5295) );
  OAI21_X4 U5998 ( .B1(n6169), .B2(n6168), .A(n6167), .ZN(n6331) );
  NAND2_X4 U5999 ( .A1(n6516), .A2(n6726), .ZN(n6367) );
  NAND2_X4 U6000 ( .A1(n4130), .A2(n4131), .ZN(n4735) );
  NAND2_X4 U6001 ( .A1(n5130), .A2(n5204), .ZN(n5209) );
  NAND2_X4 U6002 ( .A1(n5558), .A2(n5557), .ZN(n5898) );
  NAND2_X4 U6003 ( .A1(net223234), .A2(net218236), .ZN(n3810) );
  NAND2_X4 U6004 ( .A1(n3809), .A2(n3810), .ZN(net218268) );
  NAND2_X4 U6005 ( .A1(net218538), .A2(a[3]), .ZN(n3863) );
  NAND2_X4 U6006 ( .A1(n6799), .A2(n3797), .ZN(n6888) );
  INV_X4 U6007 ( .A(net213609), .ZN(net213683) );
  NAND2_X4 U6008 ( .A1(n3795), .A2(n5267), .ZN(n5396) );
  NOR2_X4 U6009 ( .A1(net216222), .A2(net216221), .ZN(n5392) );
  NAND2_X4 U6010 ( .A1(n5257), .A2(n5256), .ZN(n5391) );
  NAND2_X4 U6011 ( .A1(n5533), .A2(n5534), .ZN(n5632) );
  INV_X4 U6012 ( .A(n5535), .ZN(n5533) );
  NAND2_X2 U6013 ( .A1(net213612), .A2(net213609), .ZN(n6829) );
  NAND2_X4 U6014 ( .A1(n6612), .A2(n6667), .ZN(n6613) );
  NAND2_X4 U6015 ( .A1(n3982), .A2(net219116), .ZN(n3984) );
  NAND2_X2 U6016 ( .A1(n6486), .A2(n6485), .ZN(n3811) );
  AND2_X2 U6017 ( .A1(n6446), .A2(n6445), .ZN(n3812) );
  NOR2_X4 U6018 ( .A1(n3812), .A2(n6444), .ZN(n6448) );
  NAND2_X2 U6019 ( .A1(n6486), .A2(n6485), .ZN(n6664) );
  NAND2_X4 U6020 ( .A1(b[22]), .A2(a[1]), .ZN(n6445) );
  NAND2_X4 U6021 ( .A1(n6242), .A2(n6241), .ZN(n6409) );
  NAND2_X4 U6022 ( .A1(n6029), .A2(n6028), .ZN(n6158) );
  NAND2_X4 U6023 ( .A1(n6422), .A2(n6421), .ZN(net214459) );
  NAND2_X4 U6024 ( .A1(n6372), .A2(n3783), .ZN(n6720) );
  INV_X4 U6025 ( .A(n5414), .ZN(n5412) );
  INV_X4 U6026 ( .A(n5978), .ZN(n5976) );
  INV_X2 U6027 ( .A(net214879), .ZN(net223182) );
  NAND2_X2 U6028 ( .A1(n6287), .A2(n6288), .ZN(n6270) );
  NAND3_X2 U6029 ( .A1(n5624), .A2(n5623), .A3(n5622), .ZN(n5625) );
  NAND2_X4 U6030 ( .A1(n4073), .A2(net219630), .ZN(net218220) );
  AOI21_X4 U6031 ( .B1(n5429), .B2(n5621), .A(n5562), .ZN(n5563) );
  NAND2_X4 U6032 ( .A1(n5812), .A2(n5813), .ZN(n6026) );
  INV_X4 U6033 ( .A(n6287), .ZN(n6290) );
  OAI21_X2 U6034 ( .B1(n5635), .B2(n5637), .A(n5636), .ZN(n5532) );
  NAND2_X4 U6035 ( .A1(n6209), .A2(n6208), .ZN(n6310) );
  NAND2_X4 U6036 ( .A1(n5230), .A2(n5496), .ZN(n5491) );
  NAND2_X4 U6037 ( .A1(net216436), .A2(n5229), .ZN(n5496) );
  NAND2_X4 U6038 ( .A1(n4804), .A2(n4803), .ZN(n4981) );
  INV_X4 U6039 ( .A(n6872), .ZN(n6673) );
  NAND2_X4 U6040 ( .A1(n4158), .A2(n4159), .ZN(n4827) );
  NAND3_X1 U6041 ( .A1(n7786), .A2(n7785), .A3(n7784), .ZN(n7787) );
  NAND2_X1 U6042 ( .A1(n3362), .A2(n7583), .ZN(n7584) );
  NAND3_X1 U6043 ( .A1(n7773), .A2(n7772), .A3(n7771), .ZN(n7774) );
  NAND2_X1 U6044 ( .A1(n7588), .A2(n7773), .ZN(n7769) );
  NAND2_X1 U6045 ( .A1(n7587), .A2(n7586), .ZN(n7588) );
  OAI211_X2 U6046 ( .C1(net212672), .C2(net212673), .A(net212674), .B(
        net212061), .ZN(net212660) );
  XNOR2_X2 U6047 ( .A(net213755), .B(net213756), .ZN(net213751) );
  NAND2_X4 U6048 ( .A1(n3817), .A2(net213759), .ZN(net213442) );
  NAND2_X2 U6049 ( .A1(n3816), .A2(net213758), .ZN(net213201) );
  INV_X4 U6050 ( .A(net213759), .ZN(n3816) );
  XNOR2_X2 U6051 ( .A(net212114), .B(n3818), .ZN(net212113) );
  XNOR2_X2 U6052 ( .A(net212116), .B(n3819), .ZN(n3818) );
  XNOR2_X2 U6053 ( .A(n3820), .B(n3821), .ZN(n3819) );
  XNOR2_X2 U6054 ( .A(n3822), .B(n3823), .ZN(n3820) );
  NAND3_X2 U6055 ( .A1(net212125), .A2(net212126), .A3(net212127), .ZN(n3823)
         );
  INV_X4 U6056 ( .A(net212128), .ZN(net212127) );
  XNOR2_X2 U6057 ( .A(net212129), .B(n3824), .ZN(n3822) );
  XNOR2_X2 U6058 ( .A(n3825), .B(n3826), .ZN(n3824) );
  NOR2_X1 U6059 ( .A1(n3832), .A2(net212134), .ZN(n3826) );
  XNOR2_X1 U6060 ( .A(net212447), .B(net212140), .ZN(n3832) );
  XNOR2_X2 U6061 ( .A(n3827), .B(n3828), .ZN(n3825) );
  INV_X4 U6062 ( .A(net212140), .ZN(n3829) );
  XNOR2_X2 U6063 ( .A(net212141), .B(n3830), .ZN(n3827) );
  XNOR2_X2 U6064 ( .A(net212143), .B(n3831), .ZN(n3830) );
  NAND2_X1 U6065 ( .A1(net212145), .A2(net219468), .ZN(n3831) );
  CLKBUF_X3 U6066 ( .A(net212146), .Z(net219468) );
  INV_X4 U6067 ( .A(net215590), .ZN(n3833) );
  OAI21_X4 U6068 ( .B1(n3834), .B2(n3835), .A(net215782), .ZN(net215344) );
  INV_X4 U6069 ( .A(net215786), .ZN(n3835) );
  INV_X4 U6070 ( .A(n3836), .ZN(n3834) );
  NAND2_X2 U6071 ( .A1(net215790), .A2(net215791), .ZN(n3836) );
  NAND2_X2 U6072 ( .A1(net215584), .A2(net215585), .ZN(net215346) );
  XNOR2_X2 U6073 ( .A(net215586), .B(net215798), .ZN(net215585) );
  INV_X4 U6074 ( .A(net215799), .ZN(net215584) );
  NAND2_X4 U6075 ( .A1(net218148), .A2(net218146), .ZN(net217291) );
  INV_X4 U6076 ( .A(net218234), .ZN(net218148) );
  NAND3_X2 U6077 ( .A1(n3839), .A2(net218148), .A3(net218257), .ZN(net218244)
         );
  INV_X4 U6078 ( .A(net218240), .ZN(net218147) );
  NAND2_X4 U6079 ( .A1(net218145), .A2(net218146), .ZN(net217293) );
  INV_X8 U6080 ( .A(net218241), .ZN(net218145) );
  NAND2_X4 U6081 ( .A1(n3837), .A2(net218210), .ZN(net217294) );
  XNOR2_X2 U6082 ( .A(net218214), .B(n3206), .ZN(n3838) );
  XNOR2_X2 U6083 ( .A(net218214), .B(n3206), .ZN(net219965) );
  INV_X4 U6084 ( .A(net218146), .ZN(net218235) );
  NAND3_X1 U6085 ( .A1(net218241), .A2(net218234), .A3(net218240), .ZN(
        net218245) );
  AOI21_X2 U6086 ( .B1(net218233), .B2(net218234), .A(net218235), .ZN(
        net218206) );
  INV_X4 U6087 ( .A(net218210), .ZN(net218212) );
  XNOR2_X2 U6088 ( .A(n3847), .B(n3848), .ZN(n3846) );
  NAND2_X4 U6089 ( .A1(n3846), .A2(net214334), .ZN(net213553) );
  INV_X4 U6090 ( .A(n3846), .ZN(net214332) );
  OAI21_X4 U6091 ( .B1(n3841), .B2(n3842), .A(n3843), .ZN(net213867) );
  INV_X2 U6092 ( .A(net214338), .ZN(n3850) );
  NAND2_X2 U6093 ( .A1(n3849), .A2(net214338), .ZN(n3840) );
  INV_X2 U6094 ( .A(n3840), .ZN(net213864) );
  NAND2_X2 U6095 ( .A1(net213867), .A2(n3840), .ZN(net214038) );
  INV_X4 U6096 ( .A(net214339), .ZN(n3849) );
  OAI21_X4 U6097 ( .B1(n3851), .B2(n3852), .A(n3853), .ZN(n3844) );
  INV_X4 U6098 ( .A(n3844), .ZN(n3842) );
  INV_X4 U6099 ( .A(net214433), .ZN(n3852) );
  INV_X4 U6100 ( .A(n3845), .ZN(n3841) );
  INV_X4 U6101 ( .A(net219859), .ZN(n3854) );
  INV_X4 U6102 ( .A(net214612), .ZN(n3855) );
  NAND2_X2 U6103 ( .A1(net214433), .A2(net214434), .ZN(net214610) );
  NAND2_X2 U6104 ( .A1(net214434), .A2(net214705), .ZN(net214603) );
  NAND2_X2 U6105 ( .A1(net214612), .A2(net219859), .ZN(n3853) );
  XNOR2_X2 U6106 ( .A(net218144), .B(net218110), .ZN(net218114) );
  INV_X4 U6107 ( .A(net212688), .ZN(net212687) );
  XNOR2_X2 U6108 ( .A(n3858), .B(net216096), .ZN(n3857) );
  INV_X2 U6109 ( .A(n3785), .ZN(net216196) );
  NAND3_X4 U6110 ( .A1(n3857), .A2(net216203), .A3(n3163), .ZN(net216092) );
  INV_X1 U6111 ( .A(n3856), .ZN(n3862) );
  INV_X4 U6112 ( .A(net216022), .ZN(n3856) );
  NAND2_X4 U6113 ( .A1(net216020), .A2(n3856), .ZN(net215812) );
  INV_X1 U6114 ( .A(net216019), .ZN(net216206) );
  NAND2_X4 U6115 ( .A1(b[8]), .A2(a[8]), .ZN(net216097) );
  NAND2_X2 U6116 ( .A1(n3859), .A2(net216213), .ZN(net215813) );
  INV_X4 U6117 ( .A(net216211), .ZN(n3859) );
  INV_X4 U6118 ( .A(n3863), .ZN(net218236) );
  NAND2_X2 U6119 ( .A1(net217795), .A2(n3863), .ZN(net217427) );
  OAI22_X2 U6120 ( .A1(n3863), .A2(net218600), .B1(net218640), .B2(net217427), 
        .ZN(net217771) );
  AOI21_X4 U6121 ( .B1(n3864), .B2(net214619), .A(net214620), .ZN(net214617)
         );
  NAND2_X2 U6122 ( .A1(n3869), .A2(net215127), .ZN(n3866) );
  NAND2_X4 U6123 ( .A1(n3866), .A2(n3867), .ZN(net215124) );
  INV_X4 U6124 ( .A(net215126), .ZN(n3869) );
  NAND2_X4 U6125 ( .A1(n3868), .A2(net215126), .ZN(n3867) );
  NOR2_X4 U6126 ( .A1(n3593), .A2(n4933), .ZN(n3870) );
  INV_X4 U6127 ( .A(n3870), .ZN(n5289) );
  NAND2_X1 U6128 ( .A1(b[11]), .A2(a[1]), .ZN(n4933) );
  XOR2_X2 U6129 ( .A(n6230), .B(n6302), .Z(n3871) );
  NAND2_X4 U6130 ( .A1(n6303), .A2(n6499), .ZN(n6230) );
  XNOR2_X2 U6131 ( .A(n5567), .B(n5716), .ZN(n3872) );
  INV_X4 U6132 ( .A(net220496), .ZN(net214376) );
  NAND2_X4 U6133 ( .A1(n5896), .A2(n5898), .ZN(n5705) );
  NAND2_X4 U6134 ( .A1(n5900), .A2(n5897), .ZN(n5704) );
  NAND2_X2 U6135 ( .A1(net214834), .A2(net215468), .ZN(n5853) );
  XNOR2_X2 U6136 ( .A(n7267), .B(net213138), .ZN(n7134) );
  XNOR2_X2 U6137 ( .A(n5419), .B(n5418), .ZN(n3875) );
  AOI21_X4 U6138 ( .B1(n5425), .B2(n3886), .A(n5417), .ZN(n5418) );
  XNOR2_X1 U6139 ( .A(n6051), .B(n6049), .ZN(n3963) );
  XNOR2_X1 U6140 ( .A(n7416), .B(n7297), .ZN(n3876) );
  NAND2_X4 U6141 ( .A1(n7417), .A2(n7415), .ZN(n7297) );
  XNOR2_X2 U6142 ( .A(n5561), .B(n5563), .ZN(n3877) );
  INV_X4 U6143 ( .A(n3877), .ZN(n5565) );
  XNOR2_X2 U6144 ( .A(n3423), .B(net212656), .ZN(n7109) );
  XNOR2_X2 U6145 ( .A(n3872), .B(n3932), .ZN(net220410) );
  NAND3_X2 U6146 ( .A1(a[3]), .A2(a[2]), .A3(n4674), .ZN(n4027) );
  INV_X16 U6147 ( .A(a[3]), .ZN(net218470) );
  CLKBUF_X3 U6148 ( .A(net218273), .Z(net220397) );
  NAND2_X4 U6149 ( .A1(b[1]), .A2(b[0]), .ZN(net220396) );
  NAND2_X4 U6150 ( .A1(a[0]), .A2(a[1]), .ZN(net220394) );
  XNOR2_X2 U6151 ( .A(n5960), .B(n5959), .ZN(net220385) );
  NAND2_X1 U6152 ( .A1(n4358), .A2(net218566), .ZN(n4361) );
  NOR2_X2 U6153 ( .A1(a[1]), .A2(net218566), .ZN(n4598) );
  INV_X4 U6154 ( .A(net218566), .ZN(net218562) );
  NAND3_X2 U6155 ( .A1(n5949), .A2(n5948), .A3(n5675), .ZN(n5950) );
  NOR2_X4 U6156 ( .A1(n3893), .A2(n3353), .ZN(n3878) );
  INV_X4 U6157 ( .A(net220293), .ZN(net216008) );
  NAND2_X4 U6158 ( .A1(n5650), .A2(n3197), .ZN(n5506) );
  NAND2_X4 U6159 ( .A1(n5664), .A2(n5665), .ZN(n5796) );
  XNOR2_X2 U6160 ( .A(n7583), .B(n3362), .ZN(n3879) );
  INV_X4 U6161 ( .A(n3879), .ZN(n7547) );
  OAI21_X1 U6162 ( .B1(n7555), .B2(net220079), .A(n7554), .ZN(n7556) );
  INV_X4 U6163 ( .A(net219673), .ZN(net219674) );
  XNOR2_X2 U6164 ( .A(n5693), .B(net215770), .ZN(n3884) );
  INV_X2 U6165 ( .A(n5550), .ZN(n3885) );
  INV_X4 U6166 ( .A(n3885), .ZN(n3886) );
  NAND3_X1 U6167 ( .A1(a[24]), .A2(n7134), .A3(b[4]), .ZN(n3887) );
  XNOR2_X2 U6168 ( .A(net215124), .B(net215122), .ZN(n3950) );
  INV_X4 U6169 ( .A(net215124), .ZN(net215121) );
  XNOR2_X2 U6170 ( .A(n5297), .B(n5342), .ZN(n3888) );
  XNOR2_X2 U6171 ( .A(n5545), .B(n5537), .ZN(n3889) );
  NAND2_X4 U6172 ( .A1(n5632), .A2(net215674), .ZN(n5537) );
  NAND2_X4 U6173 ( .A1(n6094), .A2(n6093), .ZN(n6295) );
  OAI21_X4 U6174 ( .B1(n3976), .B2(n6092), .A(n6255), .ZN(n6094) );
  NAND2_X4 U6175 ( .A1(n6876), .A2(n6873), .ZN(n6614) );
  NAND2_X4 U6176 ( .A1(net213141), .A2(n7023), .ZN(net213140) );
  NAND2_X2 U6177 ( .A1(net215786), .A2(n5688), .ZN(net215783) );
  NAND2_X4 U6178 ( .A1(b[18]), .A2(a[5]), .ZN(net214549) );
  NAND2_X4 U6179 ( .A1(n4718), .A2(n4719), .ZN(n4888) );
  XNOR2_X2 U6180 ( .A(n6098), .B(n6292), .ZN(n6121) );
  INV_X4 U6181 ( .A(n6292), .ZN(n6296) );
  NAND3_X4 U6182 ( .A1(a[0]), .A2(n6097), .A3(b[20]), .ZN(n6292) );
  NOR2_X4 U6183 ( .A1(n6971), .A2(n3370), .ZN(n3890) );
  INV_X4 U6184 ( .A(n3890), .ZN(n7010) );
  NAND2_X4 U6185 ( .A1(net214732), .A2(net214731), .ZN(n6300) );
  NAND2_X4 U6186 ( .A1(n5525), .A2(n5523), .ZN(n5277) );
  INV_X4 U6187 ( .A(n5639), .ZN(n5641) );
  NOR2_X4 U6188 ( .A1(n3891), .A2(n3361), .ZN(net220099) );
  XNOR2_X2 U6189 ( .A(net213380), .B(net213381), .ZN(n3891) );
  INV_X2 U6190 ( .A(n6603), .ZN(n6601) );
  NAND2_X4 U6191 ( .A1(n5275), .A2(n5276), .ZN(n5523) );
  XOR2_X2 U6192 ( .A(n4750), .B(n4749), .Z(n3892) );
  XNOR2_X2 U6193 ( .A(n6704), .B(n6582), .ZN(n3893) );
  XNOR2_X2 U6194 ( .A(n7544), .B(n7367), .ZN(n3894) );
  XNOR2_X2 U6195 ( .A(n5411), .B(n5410), .ZN(n3895) );
  NAND2_X4 U6196 ( .A1(n5633), .A2(n5629), .ZN(n5410) );
  XOR2_X1 U6197 ( .A(n7549), .B(n7783), .Z(n3896) );
  NAND2_X4 U6198 ( .A1(n7786), .A2(n7785), .ZN(n7549) );
  NAND2_X4 U6199 ( .A1(a[10]), .A2(b[20]), .ZN(n7783) );
  NAND2_X4 U6200 ( .A1(n7568), .A2(net212126), .ZN(net212433) );
  XNOR2_X2 U6201 ( .A(n5546), .B(n5545), .ZN(n3897) );
  XNOR2_X2 U6202 ( .A(n7367), .B(n3882), .ZN(n3898) );
  INV_X1 U6203 ( .A(n4328), .ZN(n4329) );
  INV_X4 U6204 ( .A(n7027), .ZN(n7028) );
  INV_X2 U6205 ( .A(n5891), .ZN(n5847) );
  XNOR2_X2 U6206 ( .A(n5272), .B(n5271), .ZN(n3899) );
  INV_X2 U6207 ( .A(net212495), .ZN(net212493) );
  BUF_X4 U6208 ( .A(n7777), .Z(n3900) );
  NAND3_X2 U6209 ( .A1(b[24]), .A2(a[0]), .A3(n6840), .ZN(n6868) );
  AOI211_X2 U6210 ( .C1(n6641), .C2(n6840), .A(n6640), .B(n6639), .ZN(n6658)
         );
  OAI211_X1 U6211 ( .C1(n6840), .C2(n3991), .A(net218610), .B(n3414), .ZN(
        n6629) );
  NAND2_X4 U6212 ( .A1(n3593), .A2(n4933), .ZN(n5290) );
  XNOR2_X2 U6213 ( .A(n7323), .B(n7322), .ZN(n3901) );
  NAND2_X4 U6214 ( .A1(n7491), .A2(n7490), .ZN(n7322) );
  NAND2_X2 U6215 ( .A1(n4022), .A2(n3916), .ZN(net218322) );
  NAND2_X4 U6216 ( .A1(n4024), .A2(n4023), .ZN(net218321) );
  INV_X2 U6217 ( .A(net218143), .ZN(net218142) );
  AOI21_X2 U6218 ( .B1(n4106), .B2(net217242), .A(net218142), .ZN(net218140)
         );
  XNOR2_X2 U6219 ( .A(n6243), .B(n6245), .ZN(n3902) );
  XNOR2_X2 U6220 ( .A(n5018), .B(n5022), .ZN(n3903) );
  INV_X4 U6221 ( .A(n3903), .ZN(n5024) );
  NAND2_X2 U6222 ( .A1(n5213), .A2(n5076), .ZN(n5018) );
  XNOR2_X2 U6223 ( .A(n3969), .B(n4032), .ZN(n4034) );
  INV_X2 U6224 ( .A(n4033), .ZN(n3969) );
  OAI21_X1 U6225 ( .B1(n7458), .B2(n7457), .A(n7456), .ZN(n7460) );
  OAI21_X4 U6226 ( .B1(n3938), .B2(n3304), .A(n7262), .ZN(n7263) );
  NAND3_X1 U6227 ( .A1(n5890), .A2(n5891), .A3(n5892), .ZN(n5893) );
  INV_X1 U6228 ( .A(n5845), .ZN(n5615) );
  OAI21_X2 U6229 ( .B1(n3970), .B2(n5028), .A(n5141), .ZN(n5030) );
  NAND2_X4 U6230 ( .A1(n6159), .A2(n6320), .ZN(n6065) );
  NAND2_X2 U6231 ( .A1(net217075), .A2(n4818), .ZN(net216587) );
  XNOR2_X2 U6232 ( .A(n6072), .B(n6071), .ZN(n3904) );
  NAND2_X4 U6233 ( .A1(n6376), .A2(n6377), .ZN(n6715) );
  NAND2_X2 U6234 ( .A1(net213604), .A2(net213605), .ZN(n6943) );
  INV_X2 U6235 ( .A(n6319), .ZN(n3905) );
  INV_X2 U6236 ( .A(n6315), .ZN(n6319) );
  NAND2_X4 U6237 ( .A1(n6790), .A2(n6791), .ZN(n6897) );
  NAND2_X4 U6238 ( .A1(n6154), .A2(n6315), .ZN(n6071) );
  NAND2_X4 U6239 ( .A1(n3595), .A2(n5835), .ZN(n3906) );
  INV_X2 U6240 ( .A(n6775), .ZN(n6773) );
  XNOR2_X2 U6241 ( .A(net215072), .B(net215073), .ZN(n3907) );
  XNOR2_X2 U6242 ( .A(n6606), .B(n6605), .ZN(n3911) );
  NAND2_X4 U6243 ( .A1(n6678), .A2(n6939), .ZN(n6605) );
  CLKBUF_X2 U6244 ( .A(n5117), .Z(n3912) );
  NAND2_X4 U6245 ( .A1(n6593), .A2(n6594), .ZN(net213988) );
  XNOR2_X2 U6246 ( .A(net212470), .B(n7370), .ZN(n3913) );
  NAND2_X4 U6247 ( .A1(n7551), .A2(n7550), .ZN(n7370) );
  NAND2_X2 U6248 ( .A1(net216928), .A2(net216927), .ZN(net216844) );
  INV_X2 U6249 ( .A(n3219), .ZN(net219938) );
  BUF_X4 U6250 ( .A(net214785), .Z(net219931) );
  XNOR2_X2 U6251 ( .A(n6818), .B(net213969), .ZN(n3914) );
  XNOR2_X2 U6252 ( .A(net213692), .B(n6948), .ZN(n3915) );
  NAND2_X4 U6253 ( .A1(net214172), .A2(net214173), .ZN(n6807) );
  XNOR2_X2 U6254 ( .A(n3596), .B(n3270), .ZN(n3916) );
  AOI21_X2 U6255 ( .B1(n5193), .B2(net218574), .A(n4503), .ZN(n4709) );
  NOR2_X2 U6256 ( .A1(net218576), .A2(a[0]), .ZN(n4701) );
  NOR2_X2 U6257 ( .A1(n7889), .A2(net217759), .ZN(n4333) );
  NOR2_X2 U6258 ( .A1(net218484), .A2(net217759), .ZN(n4311) );
  NOR3_X2 U6259 ( .A1(n4300), .A2(n4299), .A3(n4298), .ZN(n4301) );
  NAND2_X2 U6260 ( .A1(n6950), .A2(n6949), .ZN(net219874) );
  XNOR2_X2 U6261 ( .A(n6243), .B(n6245), .ZN(n3917) );
  NAND2_X1 U6262 ( .A1(b[5]), .A2(a[7]), .ZN(net216934) );
  NAND2_X2 U6263 ( .A1(n6779), .A2(n6780), .ZN(net213764) );
  INV_X2 U6264 ( .A(n5079), .ZN(n5010) );
  NAND2_X2 U6265 ( .A1(n5215), .A2(n5084), .ZN(n5125) );
  XNOR2_X2 U6266 ( .A(n6378), .B(net214617), .ZN(net219859) );
  INV_X2 U6267 ( .A(n6063), .ZN(n6061) );
  NAND2_X2 U6268 ( .A1(n6410), .A2(n6409), .ZN(n6243) );
  OAI21_X2 U6269 ( .B1(n6719), .B2(n6718), .A(n6717), .ZN(n6900) );
  NAND2_X2 U6270 ( .A1(n6717), .A2(n6901), .ZN(n6572) );
  INV_X1 U6271 ( .A(n6506), .ZN(n6226) );
  CLKBUF_X2 U6272 ( .A(n6691), .Z(n3918) );
  NAND2_X4 U6273 ( .A1(n3892), .A2(n4751), .ZN(n4834) );
  NAND2_X4 U6274 ( .A1(n7543), .A2(n7541), .ZN(n7367) );
  NAND2_X4 U6275 ( .A1(n7364), .A2(n7365), .ZN(n7543) );
  NAND2_X4 U6276 ( .A1(net213702), .A2(net213703), .ZN(net213244) );
  NAND2_X4 U6277 ( .A1(n6814), .A2(n3954), .ZN(net213703) );
  XNOR2_X1 U6278 ( .A(n7537), .B(n7770), .ZN(n3919) );
  NAND2_X4 U6279 ( .A1(n7773), .A2(n7772), .ZN(n7537) );
  OAI21_X1 U6280 ( .B1(n7529), .B2(n7528), .A(n7527), .ZN(n7765) );
  INV_X1 U6281 ( .A(n7525), .ZN(n7529) );
  INV_X1 U6282 ( .A(n5303), .ZN(n5300) );
  INV_X4 U6283 ( .A(net219770), .ZN(net219771) );
  XNOR2_X2 U6284 ( .A(n5970), .B(net215298), .ZN(n3920) );
  OAI21_X4 U6285 ( .B1(n5888), .B2(n5887), .A(n6015), .ZN(n5970) );
  XNOR2_X2 U6286 ( .A(n6403), .B(n6404), .ZN(n3921) );
  NOR2_X4 U6287 ( .A1(n5469), .A2(n5470), .ZN(n5284) );
  INV_X2 U6288 ( .A(n5008), .ZN(n4880) );
  INV_X8 U6289 ( .A(n4730), .ZN(n4796) );
  XNOR2_X2 U6290 ( .A(net220079), .B(n7374), .ZN(n3923) );
  XNOR2_X2 U6291 ( .A(n7421), .B(n7422), .ZN(n3925) );
  INV_X4 U6292 ( .A(n3925), .ZN(n7295) );
  XNOR2_X2 U6293 ( .A(n5699), .B(n5698), .ZN(n3927) );
  NAND2_X4 U6294 ( .A1(n5907), .A2(n5903), .ZN(n5698) );
  XNOR2_X2 U6295 ( .A(net212483), .B(n7363), .ZN(n3928) );
  INV_X4 U6296 ( .A(net212485), .ZN(net212483) );
  NAND2_X4 U6297 ( .A1(n6665), .A2(n3811), .ZN(n6620) );
  NAND2_X2 U6298 ( .A1(n6941), .A2(net213607), .ZN(n6942) );
  CLKBUF_X3 U6299 ( .A(n5943), .Z(n3930) );
  NAND2_X4 U6300 ( .A1(net212137), .A2(net212138), .ZN(net212447) );
  NAND2_X1 U6301 ( .A1(n6725), .A2(n3203), .ZN(n6766) );
  NAND2_X4 U6302 ( .A1(net215786), .A2(net215782), .ZN(n5526) );
  OAI211_X2 U6303 ( .C1(n3969), .C2(n4010), .A(n4009), .B(n4119), .ZN(n4015)
         );
  OAI21_X2 U6304 ( .B1(n7520), .B2(n7519), .A(n7518), .ZN(n7521) );
  NAND2_X4 U6305 ( .A1(n7347), .A2(n7346), .ZN(n7518) );
  INV_X2 U6306 ( .A(net219678), .ZN(net219679) );
  NAND2_X4 U6307 ( .A1(n7539), .A2(n7538), .ZN(n7363) );
  NAND2_X4 U6308 ( .A1(net214853), .A2(net223422), .ZN(n6302) );
  OAI21_X2 U6309 ( .B1(n7486), .B2(n7485), .A(n7484), .ZN(n7487) );
  INV_X4 U6310 ( .A(net212656), .ZN(net212653) );
  NAND2_X4 U6311 ( .A1(n6698), .A2(n6885), .ZN(n6802) );
  NAND2_X4 U6312 ( .A1(a[2]), .A2(a[1]), .ZN(n4018) );
  XNOR2_X2 U6313 ( .A(n7485), .B(n7313), .ZN(n3933) );
  OAI21_X2 U6314 ( .B1(n7258), .B2(net212886), .A(n7257), .ZN(n7483) );
  NAND2_X2 U6315 ( .A1(n6413), .A2(n6414), .ZN(n6687) );
  NAND2_X4 U6316 ( .A1(n6947), .A2(n6946), .ZN(net213608) );
  INV_X2 U6317 ( .A(n6945), .ZN(n6947) );
  INV_X2 U6318 ( .A(n7521), .ZN(n7523) );
  NAND2_X4 U6319 ( .A1(n7522), .A2(n7521), .ZN(n7761) );
  INV_X1 U6320 ( .A(n7550), .ZN(n7552) );
  INV_X2 U6321 ( .A(net218224), .ZN(net219630) );
  INV_X4 U6322 ( .A(n4905), .ZN(n3934) );
  INV_X4 U6323 ( .A(n4142), .ZN(n3935) );
  INV_X4 U6324 ( .A(n5127), .ZN(n3936) );
  NAND2_X4 U6325 ( .A1(n4120), .A2(n4119), .ZN(n4121) );
  AOI21_X1 U6326 ( .B1(n6271), .B2(net212094), .A(n6276), .ZN(n6275) );
  INV_X1 U6327 ( .A(n6676), .ZN(n3937) );
  INV_X4 U6328 ( .A(net219569), .ZN(net218079) );
  NAND2_X2 U6329 ( .A1(net217142), .A2(net218084), .ZN(net217275) );
  NAND2_X2 U6330 ( .A1(n6965), .A2(n6966), .ZN(net219561) );
  NAND2_X2 U6331 ( .A1(n6965), .A2(n6966), .ZN(n7112) );
  INV_X2 U6332 ( .A(net219556), .ZN(net219557) );
  NOR2_X4 U6333 ( .A1(n6879), .A2(n6880), .ZN(n6882) );
  NAND2_X4 U6334 ( .A1(n7292), .A2(n7291), .ZN(n7141) );
  NAND3_X4 U6335 ( .A1(net218267), .A2(net218266), .A3(net218257), .ZN(
        net218241) );
  INV_X2 U6336 ( .A(n7375), .ZN(n7207) );
  OAI221_X1 U6337 ( .B1(n7206), .B2(net218600), .C1(n7375), .C2(n7888), .A(
        net218610), .ZN(n7210) );
  NAND2_X2 U6338 ( .A1(net213367), .A2(n7027), .ZN(n7102) );
  XNOR2_X2 U6339 ( .A(n5008), .B(n3350), .ZN(n4832) );
  NAND2_X2 U6340 ( .A1(n4999), .A2(n3943), .ZN(n5086) );
  XOR2_X2 U6341 ( .A(n7174), .B(n7173), .Z(n3939) );
  INV_X2 U6342 ( .A(n7245), .ZN(n7180) );
  XNOR2_X2 U6343 ( .A(net214840), .B(n6239), .ZN(n3940) );
  NAND2_X4 U6344 ( .A1(n5214), .A2(n5213), .ZN(n5349) );
  OAI21_X4 U6345 ( .B1(n5802), .B2(n5942), .A(n5949), .ZN(n5809) );
  AOI21_X2 U6346 ( .B1(n4844), .B2(n4843), .A(n4842), .ZN(n4846) );
  NAND2_X4 U6347 ( .A1(n5682), .A2(n5683), .ZN(net215363) );
  XNOR2_X2 U6348 ( .A(n5248), .B(n5247), .ZN(n3942) );
  NAND2_X4 U6349 ( .A1(n7109), .A2(n7110), .ZN(n7233) );
  NAND2_X4 U6350 ( .A1(n6700), .A2(n6699), .ZN(n6704) );
  XNOR2_X2 U6351 ( .A(n5241), .B(n5242), .ZN(n3943) );
  INV_X4 U6352 ( .A(n3943), .ZN(n5000) );
  NAND2_X4 U6353 ( .A1(n5001), .A2(n5000), .ZN(n5222) );
  INV_X4 U6354 ( .A(n3944), .ZN(n3945) );
  OAI21_X4 U6355 ( .B1(n3303), .B2(n3963), .A(n6162), .ZN(n6030) );
  NAND2_X4 U6356 ( .A1(net214538), .A2(n6423), .ZN(n6681) );
  XNOR2_X2 U6357 ( .A(n5516), .B(n5515), .ZN(n3946) );
  NAND2_X4 U6358 ( .A1(n6960), .A2(n6961), .ZN(n7013) );
  NAND2_X4 U6359 ( .A1(n6958), .A2(n6959), .ZN(n6961) );
  INV_X1 U6360 ( .A(n5638), .ZN(n5642) );
  INV_X8 U6361 ( .A(n5889), .ZN(n5770) );
  XNOR2_X1 U6362 ( .A(n7455), .B(n7457), .ZN(n3948) );
  XNOR2_X2 U6363 ( .A(n5681), .B(n5680), .ZN(n3949) );
  NAND2_X4 U6364 ( .A1(n5776), .A2(n5773), .ZN(n5680) );
  XNOR2_X2 U6365 ( .A(n6690), .B(n6590), .ZN(n3951) );
  XNOR2_X2 U6366 ( .A(n6392), .B(n6391), .ZN(n3952) );
  NAND2_X4 U6367 ( .A1(n6504), .A2(n6501), .ZN(n6391) );
  INV_X4 U6368 ( .A(net213612), .ZN(net213684) );
  NAND3_X2 U6369 ( .A1(n3195), .A2(net213612), .A3(n6956), .ZN(n6871) );
  INV_X2 U6370 ( .A(net212451), .ZN(net212448) );
  NAND2_X2 U6371 ( .A1(n6792), .A2(n3977), .ZN(n6895) );
  NAND2_X4 U6372 ( .A1(n5020), .A2(n5019), .ZN(n4840) );
  XNOR2_X2 U6373 ( .A(n6813), .B(n6812), .ZN(n3954) );
  NAND2_X4 U6374 ( .A1(n6686), .A2(n3421), .ZN(n6813) );
  XNOR2_X2 U6375 ( .A(n3955), .B(n3587), .ZN(n4306) );
  AND2_X2 U6376 ( .A1(net218276), .A2(net220153), .ZN(n3955) );
  NAND2_X2 U6377 ( .A1(n6690), .A2(n6689), .ZN(n6692) );
  XNOR2_X2 U6378 ( .A(net215059), .B(n6252), .ZN(n3956) );
  NAND2_X2 U6379 ( .A1(n5112), .A2(n5111), .ZN(n5115) );
  INV_X4 U6380 ( .A(n5389), .ZN(n5387) );
  XNOR2_X1 U6381 ( .A(n7167), .B(n7166), .ZN(n3957) );
  OAI21_X4 U6382 ( .B1(n5770), .B2(n5720), .A(net215477), .ZN(n5721) );
  XNOR2_X2 U6383 ( .A(n5526), .B(n5688), .ZN(n3959) );
  XNOR2_X2 U6384 ( .A(n3961), .B(n5757), .ZN(n3960) );
  AND2_X2 U6385 ( .A1(n5758), .A2(n5862), .ZN(n3961) );
  XNOR2_X2 U6386 ( .A(n5508), .B(n5645), .ZN(n3962) );
  OAI21_X2 U6387 ( .B1(net211946), .B2(n7890), .A(b[30]), .ZN(net211939) );
  NAND2_X4 U6388 ( .A1(n3317), .A2(n6048), .ZN(n6167) );
  NAND2_X4 U6389 ( .A1(n5250), .A2(n5251), .ZN(n5352) );
  NAND2_X4 U6390 ( .A1(n6694), .A2(n6697), .ZN(n6412) );
  CLKBUF_X3 U6391 ( .A(n6685), .Z(n3967) );
  XNOR2_X2 U6392 ( .A(n4996), .B(n4995), .ZN(n3968) );
  OAI21_X4 U6393 ( .B1(n5103), .B2(n5098), .A(n5104), .ZN(n4996) );
  XNOR2_X2 U6394 ( .A(n4125), .B(n3280), .ZN(net219358) );
  NAND2_X4 U6395 ( .A1(n4118), .A2(net218093), .ZN(n4125) );
  INV_X4 U6396 ( .A(n5287), .ZN(n5294) );
  NAND2_X4 U6397 ( .A1(n5086), .A2(n5222), .ZN(net216783) );
  XNOR2_X2 U6398 ( .A(net218132), .B(net218133), .ZN(n3971) );
  XNOR2_X2 U6399 ( .A(n4721), .B(n4720), .ZN(n3972) );
  NAND2_X4 U6400 ( .A1(n4891), .A2(n4888), .ZN(n4720) );
  NAND3_X1 U6401 ( .A1(n5078), .A2(n5079), .A3(n5080), .ZN(n5081) );
  NAND2_X4 U6402 ( .A1(n5077), .A2(n5073), .ZN(n4923) );
  XNOR2_X2 U6403 ( .A(n5809), .B(n5808), .ZN(n3973) );
  XNOR2_X2 U6404 ( .A(n5405), .B(n5404), .ZN(n3974) );
  NAND2_X4 U6405 ( .A1(n5472), .A2(n5636), .ZN(n5404) );
  XNOR2_X2 U6406 ( .A(n7204), .B(n7205), .ZN(net219338) );
  XNOR2_X2 U6407 ( .A(n3956), .B(net219931), .ZN(n3976) );
  XNOR2_X2 U6408 ( .A(net214019), .B(net214020), .ZN(n3977) );
  INV_X4 U6409 ( .A(n3977), .ZN(n6791) );
  XNOR2_X2 U6410 ( .A(n4909), .B(n4908), .ZN(net219328) );
  NAND2_X4 U6411 ( .A1(n4907), .A2(n4972), .ZN(n4908) );
  NAND2_X2 U6412 ( .A1(n5219), .A2(net216283), .ZN(n5118) );
  OAI21_X1 U6413 ( .B1(n7552), .B2(net212468), .A(n7551), .ZN(n7790) );
  INV_X8 U6414 ( .A(n6151), .ZN(n6307) );
  NAND2_X4 U6415 ( .A1(n6408), .A2(n3921), .ZN(n6697) );
  NAND2_X2 U6416 ( .A1(n6500), .A2(n6499), .ZN(n6392) );
  INV_X1 U6417 ( .A(n6885), .ZN(n6887) );
  NAND2_X4 U6418 ( .A1(n6615), .A2(n6616), .ZN(n6666) );
  NAND2_X4 U6419 ( .A1(n6091), .A2(n6430), .ZN(n6255) );
  NAND2_X4 U6420 ( .A1(n7162), .A2(n7163), .ZN(n7252) );
  NAND2_X4 U6421 ( .A1(n6214), .A2(n6215), .ZN(net214619) );
  INV_X4 U6422 ( .A(n6213), .ZN(n6214) );
  NAND2_X4 U6423 ( .A1(n6405), .A2(n6406), .ZN(n6694) );
  NAND2_X4 U6424 ( .A1(n6707), .A2(n6705), .ZN(n6398) );
  NAND2_X4 U6425 ( .A1(n6663), .A2(n6662), .ZN(n6832) );
  NAND2_X4 U6426 ( .A1(n6621), .A2(n6622), .ZN(n6662) );
  NAND2_X4 U6427 ( .A1(net215204), .A2(n6022), .ZN(n6023) );
  NAND2_X4 U6428 ( .A1(n5281), .A2(n5282), .ZN(n5471) );
  INV_X4 U6429 ( .A(n3949), .ZN(n5685) );
  NAND2_X4 U6430 ( .A1(n5127), .A2(n5128), .ZN(n5521) );
  NAND2_X4 U6431 ( .A1(b[1]), .A2(b[0]), .ZN(n4017) );
  NAND2_X2 U6432 ( .A1(n5298), .A2(n3978), .ZN(n3979) );
  NAND2_X2 U6433 ( .A1(n3979), .A2(n5550), .ZN(n5622) );
  NAND2_X2 U6434 ( .A1(net215674), .A2(net215673), .ZN(n5693) );
  NAND2_X2 U6435 ( .A1(n4814), .A2(net223932), .ZN(net217082) );
  NAND2_X4 U6436 ( .A1(n5539), .A2(n5538), .ZN(n5342) );
  INV_X1 U6437 ( .A(n5773), .ZN(n5774) );
  AOI21_X1 U6438 ( .B1(n6712), .B2(n6713), .A(n6711), .ZN(n6714) );
  NAND2_X4 U6439 ( .A1(n4974), .A2(n4973), .ZN(n4975) );
  NAND2_X2 U6440 ( .A1(n6507), .A2(n6506), .ZN(n6385) );
  NAND2_X4 U6441 ( .A1(n6396), .A2(n3952), .ZN(n6705) );
  OAI21_X2 U6442 ( .B1(net214954), .B2(net214955), .A(n6152), .ZN(n6309) );
  INV_X4 U6443 ( .A(n5513), .ZN(n5511) );
  NAND2_X4 U6444 ( .A1(n6586), .A2(n6587), .ZN(n6689) );
  OAI21_X4 U6445 ( .B1(n3311), .B2(n3945), .A(n5798), .ZN(n5645) );
  NAND2_X4 U6446 ( .A1(n5827), .A2(n5826), .ZN(n5906) );
  NAND2_X4 U6447 ( .A1(n5486), .A2(n5485), .ZN(n5650) );
  NAND2_X4 U6448 ( .A1(n5670), .A2(n5671), .ZN(n5948) );
  NOR2_X1 U6449 ( .A1(net218534), .A2(net218470), .ZN(n4518) );
  OAI22_X1 U6450 ( .A1(n4173), .A2(net218470), .B1(n4294), .B2(n4295), .ZN(
        n4332) );
  XNOR2_X1 U6451 ( .A(n4173), .B(net218470), .ZN(n4294) );
  NAND2_X4 U6452 ( .A1(n5279), .A2(n5280), .ZN(n5473) );
  NAND2_X4 U6453 ( .A1(n3974), .A2(n5409), .ZN(n5629) );
  NAND3_X4 U6454 ( .A1(n4410), .A2(b[6]), .A3(a[0]), .ZN(n4151) );
  OAI21_X4 U6455 ( .B1(n3314), .B2(n3942), .A(n5480), .ZN(n5354) );
  OAI22_X4 U6456 ( .A1(n4998), .A2(n4997), .B1(n5090), .B2(n5089), .ZN(n5091)
         );
  NAND2_X4 U6457 ( .A1(n4094), .A2(n4095), .ZN(net218143) );
  INV_X2 U6458 ( .A(n4485), .ZN(n4359) );
  INV_X4 U6459 ( .A(n5386), .ZN(n3980) );
  INV_X8 U6460 ( .A(n4972), .ZN(n4973) );
  NAND2_X4 U6461 ( .A1(n5913), .A2(n5909), .ZN(n5531) );
  AOI21_X4 U6462 ( .B1(net218239), .B2(net219065), .A(net218215), .ZN(
        net218214) );
  NAND2_X4 U6463 ( .A1(n7190), .A2(n7189), .ZN(net212921) );
  NOR2_X4 U6464 ( .A1(n3902), .A2(n3981), .ZN(net219178) );
  NAND2_X4 U6465 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  INV_X8 U6466 ( .A(n5854), .ZN(n6013) );
  NAND2_X1 U6467 ( .A1(n5892), .A2(n5845), .ZN(n5717) );
  NAND2_X4 U6468 ( .A1(n5621), .A2(n5617), .ZN(n5430) );
  INV_X4 U6469 ( .A(n5401), .ZN(n5402) );
  XNOR2_X2 U6470 ( .A(n6626), .B(n6661), .ZN(n6627) );
  NAND2_X4 U6471 ( .A1(n7343), .A2(n7344), .ZN(n7516) );
  NAND2_X4 U6472 ( .A1(net213749), .A2(n6930), .ZN(net213567) );
  NAND2_X4 U6473 ( .A1(n6785), .A2(n6784), .ZN(net213562) );
  NOR2_X4 U6474 ( .A1(n3907), .A2(n3327), .ZN(net219162) );
  NAND2_X4 U6475 ( .A1(net213605), .A2(n6875), .ZN(n6823) );
  INV_X4 U6476 ( .A(n5263), .ZN(n5264) );
  NAND2_X4 U6477 ( .A1(n5855), .A2(n5856), .ZN(n5886) );
  NAND2_X4 U6478 ( .A1(net213738), .A2(n6934), .ZN(net213579) );
  NAND2_X4 U6479 ( .A1(n6574), .A2(n6575), .ZN(net214323) );
  OAI21_X4 U6480 ( .B1(net214145), .B2(n6709), .A(net214147), .ZN(n6896) );
  AOI21_X2 U6481 ( .B1(n6708), .B2(n6707), .A(n6706), .ZN(n6709) );
  NAND2_X4 U6482 ( .A1(n4744), .A2(n4745), .ZN(n4823) );
  NAND2_X4 U6483 ( .A1(n3316), .A2(n4155), .ZN(n4736) );
  NAND2_X4 U6484 ( .A1(n4076), .A2(n4091), .ZN(net218042) );
  NAND2_X4 U6485 ( .A1(n3417), .A2(n5852), .ZN(net215468) );
  NAND2_X4 U6486 ( .A1(n5902), .A2(n3989), .ZN(n5699) );
  AOI21_X4 U6487 ( .B1(n6244), .B2(n3639), .A(net214830), .ZN(n6245) );
  OAI21_X1 U6488 ( .B1(n7540), .B2(net212483), .A(n7539), .ZN(n7777) );
  OAI21_X4 U6489 ( .B1(n4880), .B2(n4879), .A(n5080), .ZN(n4916) );
  NAND2_X4 U6490 ( .A1(n6238), .A2(n6237), .ZN(n6493) );
  NAND3_X2 U6491 ( .A1(n3989), .A2(n5903), .A3(n5902), .ZN(n5905) );
  NAND2_X4 U6492 ( .A1(n4122), .A2(n4121), .ZN(net217142) );
  NAND2_X4 U6493 ( .A1(n5296), .A2(n5295), .ZN(n5539) );
  NAND2_X4 U6494 ( .A1(n4127), .A2(n4128), .ZN(n4730) );
  NAND2_X1 U6495 ( .A1(n5148), .A2(n5149), .ZN(n5034) );
  XNOR2_X1 U6496 ( .A(n4920), .B(n3922), .ZN(n4921) );
  NAND2_X4 U6497 ( .A1(n5691), .A2(net215773), .ZN(net215672) );
  NAND2_X2 U6498 ( .A1(net218143), .A2(n4096), .ZN(n4097) );
  NAND2_X2 U6499 ( .A1(n7102), .A2(net212705), .ZN(n7030) );
  NAND2_X4 U6500 ( .A1(n6962), .A2(n6961), .ZN(n7012) );
  NAND2_X2 U6501 ( .A1(net217083), .A2(n4724), .ZN(n3983) );
  NAND2_X4 U6502 ( .A1(n3984), .A2(n3983), .ZN(net217235) );
  INV_X4 U6503 ( .A(n4724), .ZN(n3982) );
  NAND2_X2 U6504 ( .A1(net218306), .A2(n4036), .ZN(n3986) );
  NAND2_X4 U6505 ( .A1(n3985), .A2(net219120), .ZN(n3987) );
  NAND2_X4 U6506 ( .A1(n3986), .A2(n3987), .ZN(n4054) );
  INV_X4 U6507 ( .A(net218306), .ZN(net219120) );
  INV_X4 U6508 ( .A(n4036), .ZN(n3985) );
  NAND2_X4 U6509 ( .A1(n6248), .A2(n6249), .ZN(n6425) );
  NAND2_X4 U6510 ( .A1(b[5]), .A2(a[5]), .ZN(net217083) );
  NAND2_X4 U6511 ( .A1(n4918), .A2(n4919), .ZN(n5073) );
  INV_X2 U6512 ( .A(n4022), .ZN(n4024) );
  NAND2_X4 U6513 ( .A1(n4885), .A2(n4794), .ZN(n4729) );
  INV_X4 U6514 ( .A(n5268), .ZN(n5270) );
  NAND2_X4 U6515 ( .A1(n5477), .A2(n5476), .ZN(n5386) );
  INV_X2 U6516 ( .A(net214536), .ZN(net214538) );
  INV_X4 U6517 ( .A(n6150), .ZN(n6082) );
  NAND2_X4 U6518 ( .A1(n6897), .A2(n6895), .ZN(n6793) );
  NAND2_X4 U6519 ( .A1(n6803), .A2(n6804), .ZN(net213577) );
  NAND2_X4 U6520 ( .A1(n4712), .A2(a[9]), .ZN(net217133) );
  NAND2_X4 U6521 ( .A1(n3303), .A2(n5941), .ZN(n6162) );
  INV_X1 U6522 ( .A(n7530), .ZN(n7532) );
  NAND2_X4 U6523 ( .A1(n7516), .A2(n7518), .ZN(n7348) );
  OAI21_X1 U6524 ( .B1(n7504), .B2(n7503), .A(n7502), .ZN(n7506) );
  INV_X2 U6525 ( .A(n7249), .ZN(n7250) );
  OAI21_X2 U6526 ( .B1(n7270), .B2(n7269), .A(n7268), .ZN(n7429) );
  NAND2_X4 U6527 ( .A1(n6304), .A2(n6303), .ZN(n6500) );
  NAND2_X4 U6528 ( .A1(n3615), .A2(net218276), .ZN(n4041) );
  NAND2_X2 U6529 ( .A1(n5983), .A2(net215275), .ZN(n6428) );
  NAND2_X1 U6530 ( .A1(n4827), .A2(n4825), .ZN(n4164) );
  OAI21_X2 U6531 ( .B1(n4740), .B2(n4739), .A(n4738), .ZN(n4742) );
  NAND2_X1 U6532 ( .A1(n4152), .A2(n4151), .ZN(n4153) );
  INV_X2 U6533 ( .A(n4134), .ZN(n4146) );
  NAND2_X4 U6534 ( .A1(n4134), .A2(n4135), .ZN(n4152) );
  NAND2_X1 U6535 ( .A1(n6295), .A2(n6293), .ZN(n6098) );
  INV_X2 U6536 ( .A(n5030), .ZN(n5031) );
  NAND2_X2 U6537 ( .A1(n4840), .A2(n4930), .ZN(n4844) );
  NAND2_X4 U6538 ( .A1(n7298), .A2(n3323), .ZN(n7412) );
  INV_X2 U6539 ( .A(n5341), .ZN(n5344) );
  INV_X4 U6540 ( .A(n4053), .ZN(n4052) );
  INV_X4 U6541 ( .A(n5224), .ZN(n5225) );
  NAND2_X4 U6542 ( .A1(n6687), .A2(n6489), .ZN(n6417) );
  OAI21_X4 U6543 ( .B1(n5940), .B2(n5939), .A(n5938), .ZN(n6049) );
  NAND2_X4 U6544 ( .A1(n3959), .A2(n5527), .ZN(n5913) );
  INV_X2 U6545 ( .A(n4057), .ZN(n4059) );
  NAND2_X4 U6546 ( .A1(n6301), .A2(n6493), .ZN(n6239) );
  INV_X4 U6547 ( .A(n5121), .ZN(n5119) );
  OAI21_X2 U6548 ( .B1(net215662), .B2(net215661), .A(n3571), .ZN(n5961) );
  NAND2_X4 U6549 ( .A1(n4808), .A2(n4809), .ZN(n4972) );
  INV_X4 U6550 ( .A(n4811), .ZN(n4808) );
  OAI21_X4 U6551 ( .B1(n5958), .B2(n5957), .A(n3931), .ZN(n6028) );
  NAND2_X4 U6552 ( .A1(n5237), .A2(n5238), .ZN(n5364) );
  NAND2_X4 U6553 ( .A1(n4897), .A2(n5104), .ZN(n5098) );
  NAND2_X4 U6554 ( .A1(n4722), .A2(n4723), .ZN(n4815) );
  INV_X8 U6555 ( .A(n5084), .ZN(n5218) );
  NAND2_X4 U6556 ( .A1(n5100), .A2(n5099), .ZN(n5102) );
  NAND3_X2 U6557 ( .A1(n4714), .A2(net218096), .A3(net220022), .ZN(n4118) );
  NAND2_X4 U6558 ( .A1(n4816), .A2(net217094), .ZN(net217092) );
  NAND2_X4 U6559 ( .A1(n4982), .A2(n4981), .ZN(n4904) );
  XNOR2_X2 U6560 ( .A(n4067), .B(n3909), .ZN(n4070) );
  INV_X4 U6561 ( .A(net219063), .ZN(net219036) );
  NAND2_X4 U6562 ( .A1(n5794), .A2(n3309), .ZN(n5938) );
  NAND2_X4 U6563 ( .A1(n4012), .A2(n4013), .ZN(net218269) );
  NAND2_X1 U6564 ( .A1(n3988), .A2(net218566), .ZN(n4265) );
  NAND2_X2 U6565 ( .A1(net218354), .A2(n3988), .ZN(n4028) );
  NAND2_X4 U6566 ( .A1(net218574), .A2(a[11]), .ZN(net216517) );
  NAND2_X4 U6567 ( .A1(n5373), .A2(n5374), .ZN(n5649) );
  NAND2_X4 U6568 ( .A1(n6149), .A2(n6148), .ZN(net215089) );
  NAND2_X4 U6569 ( .A1(n6591), .A2(n6592), .ZN(net213990) );
  NAND2_X4 U6570 ( .A1(n6578), .A2(n6579), .ZN(n6703) );
  INV_X2 U6571 ( .A(n6580), .ZN(n6578) );
  NOR2_X2 U6572 ( .A1(n6014), .A2(n6013), .ZN(n6016) );
  INV_X4 U6573 ( .A(net213732), .ZN(net213730) );
  NAND2_X4 U6574 ( .A1(n7146), .A2(n7145), .ZN(n7299) );
  NAND2_X4 U6575 ( .A1(n7135), .A2(n7264), .ZN(n7265) );
  NAND2_X4 U6576 ( .A1(n3936), .A2(n5126), .ZN(n5348) );
  NAND2_X4 U6577 ( .A1(n3975), .A2(n5723), .ZN(n5760) );
  NAND2_X4 U6578 ( .A1(n5530), .A2(n5529), .ZN(n5909) );
  INV_X2 U6579 ( .A(n6705), .ZN(n6706) );
  NAND2_X4 U6580 ( .A1(n6620), .A2(n6666), .ZN(n6956) );
  NAND2_X4 U6581 ( .A1(n6607), .A2(n6608), .ZN(n6876) );
  OAI21_X1 U6582 ( .B1(n7532), .B2(net212493), .A(n7531), .ZN(n7533) );
  NAND2_X4 U6583 ( .A1(n7531), .A2(n7530), .ZN(n7358) );
  NAND2_X4 U6584 ( .A1(n6689), .A2(n6691), .ZN(n6590) );
  NAND2_X4 U6585 ( .A1(n5843), .A2(n5842), .ZN(n5894) );
  NAND2_X4 U6586 ( .A1(n6881), .A2(n6877), .ZN(n6812) );
  NAND2_X4 U6587 ( .A1(n5358), .A2(n5357), .ZN(n5481) );
  NAND2_X2 U6588 ( .A1(n5481), .A2(n5480), .ZN(n5384) );
  INV_X2 U6589 ( .A(n3910), .ZN(n4358) );
  NAND2_X4 U6590 ( .A1(n5686), .A2(net215802), .ZN(net215667) );
  INV_X8 U6591 ( .A(n4982), .ZN(n4984) );
  NAND3_X4 U6592 ( .A1(n4890), .A2(n3272), .A3(n4892), .ZN(n4982) );
  NAND2_X4 U6593 ( .A1(net217077), .A2(n4817), .ZN(net216932) );
  NAND2_X4 U6594 ( .A1(n4137), .A2(n4135), .ZN(n4113) );
  INV_X2 U6595 ( .A(net213752), .ZN(net213753) );
  NAND2_X4 U6596 ( .A1(net214863), .A2(net219771), .ZN(n6222) );
  NAND2_X1 U6597 ( .A1(n4032), .A2(n4029), .ZN(n4031) );
  NAND2_X4 U6598 ( .A1(n5541), .A2(n5542), .ZN(n5630) );
  INV_X2 U6599 ( .A(net219485), .ZN(net216796) );
  NAND2_X4 U6600 ( .A1(n5387), .A2(n5388), .ZN(n5474) );
  INV_X8 U6601 ( .A(net218566), .ZN(net218560) );
  NAND2_X4 U6602 ( .A1(n3884), .A2(n5697), .ZN(n5903) );
  NAND2_X4 U6603 ( .A1(n5694), .A2(n5695), .ZN(n5907) );
  NAND2_X4 U6604 ( .A1(n6822), .A2(n6821), .ZN(n6875) );
  INV_X4 U6605 ( .A(n6820), .ZN(n6822) );
  NAND2_X4 U6606 ( .A1(n7182), .A2(n7183), .ZN(n7238) );
  NAND2_X4 U6607 ( .A1(n6217), .A2(n6218), .ZN(net214705) );
  NAND2_X4 U6608 ( .A1(net213072), .A2(n3939), .ZN(n7177) );
  NAND2_X2 U6609 ( .A1(n7112), .A2(net213375), .ZN(n6969) );
  NAND2_X4 U6610 ( .A1(n4914), .A2(n4913), .ZN(n5079) );
  NAND2_X4 U6611 ( .A1(n3172), .A2(n5706), .ZN(n5895) );
  NAND2_X4 U6612 ( .A1(n5703), .A2(n3927), .ZN(n5897) );
  INV_X4 U6613 ( .A(n6293), .ZN(n6294) );
  NAND2_X4 U6614 ( .A1(n5144), .A2(n5145), .ZN(n5200) );
  NAND2_X4 U6615 ( .A1(n3774), .A2(n4126), .ZN(n4795) );
  NAND3_X2 U6616 ( .A1(net214568), .A2(n6409), .A3(n3639), .ZN(n6411) );
  NAND3_X2 U6617 ( .A1(n5863), .A2(n5862), .A3(n5861), .ZN(net215516) );
  NAND3_X2 U6618 ( .A1(a[0]), .A2(b[18]), .A3(n3960), .ZN(n5981) );
  NAND2_X4 U6619 ( .A1(n5270), .A2(n5269), .ZN(net216200) );
  INV_X1 U6620 ( .A(n5860), .ZN(n5861) );
  NAND2_X4 U6621 ( .A1(net216200), .A2(n5396), .ZN(n5271) );
  INV_X2 U6622 ( .A(n4092), .ZN(n4066) );
  NAND2_X4 U6623 ( .A1(n4093), .A2(n4092), .ZN(net218116) );
  NAND2_X4 U6624 ( .A1(n5676), .A2(n5677), .ZN(n5776) );
  OAI221_X4 U6625 ( .B1(n5105), .B2(n5104), .C1(n5103), .C2(n5102), .A(n5101), 
        .ZN(n5231) );
  NAND2_X4 U6626 ( .A1(n5017), .A2(n5016), .ZN(n5076) );
  NAND2_X4 U6627 ( .A1(n5730), .A2(n5729), .ZN(n5758) );
  NAND2_X4 U6628 ( .A1(n5412), .A2(n5413), .ZN(n5627) );
  NAND2_X4 U6629 ( .A1(n7357), .A2(n7356), .ZN(n7530) );
  NAND2_X4 U6630 ( .A1(n7362), .A2(n7361), .ZN(n7538) );
  NOR2_X2 U6631 ( .A1(n6886), .A2(n6887), .ZN(n6889) );
  AOI21_X2 U6632 ( .B1(n4922), .B2(n5077), .A(n5021), .ZN(n5022) );
  NAND2_X2 U6633 ( .A1(net216840), .A2(n3299), .ZN(n4820) );
  NAND2_X4 U6634 ( .A1(n4084), .A2(n4083), .ZN(net218058) );
  NAND2_X4 U6635 ( .A1(n4090), .A2(n4089), .ZN(net218059) );
  NAND2_X4 U6636 ( .A1(n4037), .A2(n4045), .ZN(net218240) );
  NAND2_X4 U6637 ( .A1(n4117), .A2(n3971), .ZN(n4792) );
  NAND2_X2 U6638 ( .A1(n5014), .A2(n5015), .ZN(n5213) );
  NAND3_X2 U6639 ( .A1(n4887), .A2(n4889), .A3(n4888), .ZN(n4805) );
  NAND3_X2 U6640 ( .A1(n4887), .A2(n4888), .A3(n4889), .ZN(n4890) );
  NAND3_X2 U6641 ( .A1(n4814), .A2(net216945), .A3(net223932), .ZN(n4816) );
  NAND2_X4 U6642 ( .A1(n6393), .A2(n6394), .ZN(n6707) );
  NAND2_X4 U6643 ( .A1(n7570), .A2(n7569), .ZN(n7568) );
  NAND2_X4 U6644 ( .A1(n5406), .A2(n5407), .ZN(n5633) );
  NAND2_X4 U6645 ( .A1(n3928), .A2(n7366), .ZN(n7541) );
  NAND2_X4 U6646 ( .A1(n4839), .A2(n4838), .ZN(n4930) );
  NAND2_X4 U6647 ( .A1(n5587), .A2(n5586), .ZN(n5762) );
  NAND2_X4 U6648 ( .A1(b[1]), .A2(a[4]), .ZN(n4067) );
  OAI21_X4 U6649 ( .B1(n6025), .B2(net220385), .A(n6023), .ZN(n6155) );
  NAND2_X4 U6650 ( .A1(n4025), .A2(n4027), .ZN(n4029) );
  XNOR2_X1 U6651 ( .A(net212134), .B(n3832), .ZN(n7572) );
  XNOR2_X1 U6652 ( .A(net212145), .B(net219468), .ZN(n7576) );
  INV_X2 U6653 ( .A(net213716), .ZN(net213718) );
  NAND2_X4 U6654 ( .A1(n7352), .A2(n7351), .ZN(n7525) );
  INV_X8 U6655 ( .A(n7116), .ZN(n7273) );
  NAND2_X4 U6656 ( .A1(n6777), .A2(n6778), .ZN(net213555) );
  NAND2_X4 U6657 ( .A1(n7289), .A2(n7456), .ZN(n7457) );
  INV_X2 U6658 ( .A(n6879), .ZN(n6686) );
  NAND2_X4 U6659 ( .A1(n5140), .A2(n5139), .ZN(n5292) );
  XNOR2_X2 U6660 ( .A(n5138), .B(n3965), .ZN(n5139) );
  NAND2_X4 U6661 ( .A1(net216008), .A2(n5520), .ZN(net215782) );
  NAND2_X4 U6662 ( .A1(n5966), .A2(n5967), .ZN(net214979) );
  NAND3_X1 U6663 ( .A1(net216842), .A2(net216927), .A3(net216928), .ZN(
        net216926) );
  NAND2_X4 U6664 ( .A1(n7142), .A2(n3304), .ZN(n7262) );
  NAND2_X4 U6665 ( .A1(n5422), .A2(n5423), .ZN(n5617) );
  NAND2_X4 U6666 ( .A1(net218574), .A2(a[7]), .ZN(n4485) );
  NAND2_X2 U6667 ( .A1(n4972), .A2(n4978), .ZN(net217091) );
  NAND2_X2 U6668 ( .A1(n4811), .A2(n4810), .ZN(n4978) );
  NAND2_X4 U6669 ( .A1(n7252), .A2(n7249), .ZN(n7166) );
  NAND2_X4 U6670 ( .A1(n5265), .A2(n5264), .ZN(net216019) );
  NAND2_X2 U6671 ( .A1(n5851), .A2(n3784), .ZN(net214834) );
  NAND2_X4 U6672 ( .A1(n6017), .A2(n3282), .ZN(n5965) );
  NAND3_X2 U6673 ( .A1(n6229), .A2(n6506), .A3(n6228), .ZN(n6499) );
  NAND2_X4 U6674 ( .A1(n6222), .A2(n6223), .ZN(n6506) );
  INV_X2 U6675 ( .A(n5020), .ZN(n4838) );
  NAND3_X2 U6676 ( .A1(n6224), .A2(net219771), .A3(net214863), .ZN(n6229) );
  INV_X1 U6677 ( .A(n6625), .ZN(n6449) );
  OAI211_X4 U6678 ( .C1(n7236), .C2(n7237), .A(net212954), .B(n7235), .ZN(
        net212442) );
  NAND2_X4 U6679 ( .A1(n5356), .A2(n3806), .ZN(n5357) );
  NAND2_X4 U6680 ( .A1(n5113), .A2(n5114), .ZN(n5355) );
  OAI21_X4 U6681 ( .B1(n3958), .B2(n3313), .A(net216841), .ZN(n4791) );
  NAND2_X4 U6682 ( .A1(n4734), .A2(n3313), .ZN(net216841) );
  NOR2_X2 U6683 ( .A1(net220396), .A2(n4018), .ZN(n4020) );
  NAND3_X2 U6684 ( .A1(n6839), .A2(n6838), .A3(n6837), .ZN(net213374) );
  OAI21_X2 U6685 ( .B1(net212437), .B2(net212438), .A(net223689), .ZN(n7566)
         );
  NAND2_X4 U6686 ( .A1(n5718), .A2(n5719), .ZN(net215477) );
  INV_X2 U6687 ( .A(net212636), .ZN(net212635) );
  NAND2_X4 U6688 ( .A1(n3328), .A2(n7168), .ZN(net212636) );
  INV_X2 U6689 ( .A(n5135), .ZN(n5133) );
  NAND2_X4 U6690 ( .A1(net220293), .A2(n5519), .ZN(net215786) );
  NAND2_X4 U6691 ( .A1(n5565), .A2(n5564), .ZN(n5892) );
  NAND2_X2 U6692 ( .A1(n5222), .A2(n5223), .ZN(n5116) );
  NAND2_X4 U6693 ( .A1(net215591), .A2(net215590), .ZN(net215347) );
  NAND2_X4 U6694 ( .A1(n5420), .A2(n5421), .ZN(n5621) );
  NAND2_X2 U6695 ( .A1(net216202), .A2(n5394), .ZN(n5272) );
  NAND2_X4 U6696 ( .A1(n6811), .A2(n6810), .ZN(n6877) );
  NAND2_X4 U6697 ( .A1(n5759), .A2(n5758), .ZN(n5863) );
  NAND2_X4 U6698 ( .A1(n6827), .A2(n6828), .ZN(net213609) );
  NAND2_X4 U6699 ( .A1(n6703), .A2(n6701), .ZN(n6582) );
  NAND3_X2 U6700 ( .A1(net216001), .A2(n5525), .A3(n5524), .ZN(net215791) );
  NAND2_X4 U6701 ( .A1(n4924), .A2(n4925), .ZN(n4963) );
  NAND2_X4 U6702 ( .A1(n5303), .A2(n5302), .ZN(n5618) );
  NAND3_X2 U6703 ( .A1(n5627), .A2(n5626), .A3(n5625), .ZN(n5902) );
  NAND3_X1 U6704 ( .A1(net217242), .A2(net217240), .A3(net218114), .ZN(
        net218136) );
  NAND2_X4 U6705 ( .A1(n5121), .A2(n5122), .ZN(net216393) );
  NAND2_X4 U6706 ( .A1(n5560), .A2(n5559), .ZN(n5620) );
  NAND3_X2 U6707 ( .A1(net218244), .A2(net218245), .A3(n4064), .ZN(net218115)
         );
  NAND2_X4 U6708 ( .A1(n5403), .A2(n5402), .ZN(n5636) );
  NAND2_X4 U6709 ( .A1(net218237), .A2(net218236), .ZN(net218146) );
  NAND2_X4 U6710 ( .A1(n3917), .A2(n6247), .ZN(net214716) );
  NAND3_X2 U6711 ( .A1(n4028), .A2(n4027), .A3(n4026), .ZN(n4032) );
  NAND2_X4 U6712 ( .A1(a[3]), .A2(a[2]), .ZN(net218367) );
  NAND2_X4 U6713 ( .A1(n4103), .A2(net218166), .ZN(n4072) );
  NAND2_X1 U6714 ( .A1(a[0]), .A2(net218576), .ZN(n4700) );
  NAND2_X1 U6715 ( .A1(a[31]), .A2(net218576), .ZN(n7668) );
  NAND2_X1 U6716 ( .A1(a[30]), .A2(net218574), .ZN(n7438) );
  NAND2_X1 U6717 ( .A1(a[29]), .A2(net218574), .ZN(n7817) );
  NAND2_X1 U6718 ( .A1(a[28]), .A2(net218576), .ZN(n7217) );
  NAND2_X1 U6719 ( .A1(a[27]), .A2(net218574), .ZN(n7816) );
  NAND2_X4 U6720 ( .A1(n3923), .A2(net212738), .ZN(net212645) );
  XNOR2_X2 U6721 ( .A(n5717), .B(n3932), .ZN(n5718) );
  NAND2_X4 U6722 ( .A1(n6595), .A2(n6596), .ZN(n6682) );
  NAND2_X4 U6723 ( .A1(b[1]), .A2(a[2]), .ZN(n4006) );
  NAND2_X4 U6724 ( .A1(net218550), .A2(a[2]), .ZN(n4248) );
  NAND2_X4 U6725 ( .A1(net218536), .A2(a[2]), .ZN(n4045) );
  INV_X2 U6726 ( .A(n6884), .ZN(n6890) );
  NAND2_X4 U6727 ( .A1(n6888), .A2(n6884), .ZN(n6801) );
  NAND2_X4 U6728 ( .A1(n5431), .A2(n5432), .ZN(n5574) );
  OAI21_X4 U6729 ( .B1(n5344), .B2(n5343), .A(n5630), .ZN(n5411) );
  NAND2_X4 U6730 ( .A1(n6416), .A2(n6415), .ZN(n6489) );
  NAND2_X4 U6731 ( .A1(n6390), .A2(n6389), .ZN(n6501) );
  NAND2_X4 U6732 ( .A1(n6402), .A2(n6401), .ZN(n6495) );
  NAND3_X2 U6733 ( .A1(n5630), .A2(n5629), .A3(n5628), .ZN(n5631) );
  NAND2_X4 U6734 ( .A1(n6411), .A2(n6410), .ZN(n6693) );
  OAI21_X2 U6735 ( .B1(net214728), .B2(n6300), .A(net224078), .ZN(net214726)
         );
  NAND2_X4 U6736 ( .A1(n5976), .A2(n5977), .ZN(net215057) );
  NAND2_X4 U6737 ( .A1(n6258), .A2(n6259), .ZN(n6291) );
  NAND2_X4 U6738 ( .A1(n4929), .A2(n4841), .ZN(n4965) );
  NAND2_X4 U6739 ( .A1(n7175), .A2(net213070), .ZN(n7245) );
  NAND2_X4 U6740 ( .A1(n7527), .A2(n7525), .ZN(n7353) );
  NAND2_X4 U6741 ( .A1(n6892), .A2(n6891), .ZN(n6797) );
  OAI21_X2 U6742 ( .B1(net218273), .B2(net218308), .A(net218272), .ZN(n4036)
         );
  OAI211_X1 U6743 ( .C1(n6097), .C2(net218655), .A(net218608), .B(n3413), .ZN(
        n5991) );
  NAND2_X4 U6744 ( .A1(n4882), .A2(n4881), .ZN(net216840) );
  NAND2_X1 U6745 ( .A1(n4266), .A2(net218574), .ZN(n4449) );
  INV_X2 U6746 ( .A(n6441), .ZN(n6669) );
  NAND2_X1 U6747 ( .A1(a[13]), .A2(net218574), .ZN(net216117) );
  OAI22_X4 U6748 ( .A1(net219036), .A2(n3296), .B1(net219054), .B2(n4019), 
        .ZN(n4011) );
  NAND3_X1 U6749 ( .A1(n5617), .A2(n5618), .A3(n5616), .ZN(n5619) );
  NAND2_X4 U6750 ( .A1(n3873), .A2(n6796), .ZN(n6891) );
  NAND2_X4 U6751 ( .A1(net217817), .A2(net218558), .ZN(n5044) );
  NAND2_X4 U6752 ( .A1(n7203), .A2(n7202), .ZN(net212703) );
  OAI21_X1 U6753 ( .B1(n6262), .B2(n6292), .A(n6293), .ZN(n6263) );
  NAND2_X4 U6754 ( .A1(n3894), .A2(n7369), .ZN(n7550) );
  NAND2_X4 U6755 ( .A1(n3762), .A2(n5566), .ZN(n5845) );
  NAND2_X4 U6756 ( .A1(n6096), .A2(n6095), .ZN(n6293) );
  XNOR2_X2 U6757 ( .A(n7025), .B(net219657), .ZN(n7026) );
  NAND2_X4 U6758 ( .A1(n7102), .A2(n7103), .ZN(net212704) );
  NAND2_X4 U6759 ( .A1(net217236), .A2(net216947), .ZN(n4814) );
  NAND2_X4 U6760 ( .A1(n7028), .A2(net213364), .ZN(net212705) );
  NAND2_X4 U6761 ( .A1(n5003), .A2(n5004), .ZN(n5084) );
  NAND3_X2 U6762 ( .A1(n5621), .A2(n5620), .A3(n5619), .ZN(n5896) );
  NAND2_X4 U6763 ( .A1(net218099), .A2(net219065), .ZN(n4714) );
  OAI21_X2 U6764 ( .B1(n4008), .B2(net218352), .A(net218353), .ZN(n4010) );
  NAND2_X4 U6765 ( .A1(n5284), .A2(n3162), .ZN(n5634) );
  NAND2_X1 U6766 ( .A1(n3209), .A2(net220153), .ZN(n4038) );
  NAND2_X4 U6767 ( .A1(b[1]), .A2(b[0]), .ZN(n4019) );
  NAND2_X4 U6768 ( .A1(a[3]), .A2(b[0]), .ZN(n4005) );
  NAND2_X4 U6769 ( .A1(n3895), .A2(n5415), .ZN(n5623) );
  NAND2_X4 U6770 ( .A1(n4102), .A2(n4101), .ZN(net217242) );
  OAI21_X2 U6771 ( .B1(n3976), .B2(n6431), .A(n6429), .ZN(n6433) );
  NAND2_X4 U6772 ( .A1(net215277), .A2(n5982), .ZN(n6089) );
  NAND2_X4 U6773 ( .A1(n5700), .A2(n5701), .ZN(n5900) );
  NAND3_X2 U6774 ( .A1(n5910), .A2(n5909), .A3(n5908), .ZN(n5822) );
  NAND2_X2 U6775 ( .A1(n5636), .A2(n5637), .ZN(n5908) );
  NAND2_X4 U6776 ( .A1(n3950), .A2(n6081), .ZN(n6150) );
  NAND2_X4 U6777 ( .A1(n5507), .A2(n3311), .ZN(n5798) );
  NAND3_X2 U6778 ( .A1(n5631), .A2(n5632), .A3(n5633), .ZN(net215673) );
  INV_X8 U6779 ( .A(net216190), .ZN(net216193) );
  NAND2_X4 U6780 ( .A1(n4100), .A2(n4099), .ZN(net218043) );
  OAI21_X4 U6781 ( .B1(n3315), .B2(n3964), .A(n3210), .ZN(n5478) );
  NAND2_X1 U6782 ( .A1(n6869), .A2(net213374), .ZN(n6841) );
  NAND2_X4 U6783 ( .A1(n6870), .A2(n6869), .ZN(net213373) );
  NAND2_X1 U6784 ( .A1(n5892), .A2(n5890), .ZN(n5848) );
  NAND2_X4 U6785 ( .A1(n5892), .A2(n5845), .ZN(n5567) );
  NAND2_X4 U6786 ( .A1(n3934), .A2(n4971), .ZN(n4979) );
  NAND2_X4 U6787 ( .A1(n3773), .A2(n5821), .ZN(net215434) );
  NAND2_X4 U6788 ( .A1(n4726), .A2(n4725), .ZN(n4885) );
  NAND2_X4 U6789 ( .A1(n5093), .A2(n5092), .ZN(n5241) );
  NAND2_X4 U6790 ( .A1(n5511), .A2(n5512), .ZN(n5640) );
  NAND2_X4 U6791 ( .A1(n5117), .A2(n3312), .ZN(net216284) );
  NAND2_X4 U6792 ( .A1(n3972), .A2(n4813), .ZN(n4906) );
  NAND2_X4 U6793 ( .A1(n6817), .A2(n6816), .ZN(net213598) );
  NAND2_X4 U6794 ( .A1(n6495), .A2(n6699), .ZN(n6403) );
  NAND2_X4 U6795 ( .A1(n6024), .A2(net215206), .ZN(net215199) );
  NAND2_X4 U6796 ( .A1(n5810), .A2(n3321), .ZN(n5956) );
  INV_X2 U6797 ( .A(n5946), .ZN(n5802) );
  NAND2_X4 U6798 ( .A1(n5711), .A2(n5712), .ZN(net215478) );
  NAND2_X4 U6799 ( .A1(n5002), .A2(n3308), .ZN(net216283) );
  NAND2_X4 U6800 ( .A1(n5119), .A2(n5120), .ZN(net216219) );
  NAND2_X4 U6801 ( .A1(net217281), .A2(n4889), .ZN(n4721) );
  NAND2_X4 U6802 ( .A1(n5685), .A2(n5684), .ZN(net215663) );
  OAI21_X2 U6803 ( .B1(net216251), .B2(n5495), .A(n5494), .ZN(n5371) );
  NAND2_X4 U6804 ( .A1(n3204), .A2(n5673), .ZN(n5943) );
  NAND2_X4 U6805 ( .A1(n3914), .A2(n6819), .ZN(net213605) );
  NAND2_X4 U6806 ( .A1(n5707), .A2(n5708), .ZN(n5891) );
  NAND2_X4 U6807 ( .A1(n5627), .A2(n5623), .ZN(n5416) );
  NAND3_X2 U6808 ( .A1(n4977), .A2(n4978), .A3(net216819), .ZN(n4907) );
  NAND2_X4 U6809 ( .A1(n4815), .A2(n4906), .ZN(net216941) );
  NOR2_X4 U6810 ( .A1(net215662), .A2(net215661), .ZN(net215805) );
  NAND2_X4 U6811 ( .A1(net217118), .A2(n4798), .ZN(n4986) );
  NAND2_X4 U6812 ( .A1(n4715), .A2(n4716), .ZN(n4891) );
  NAND2_X4 U6813 ( .A1(n4048), .A2(n4047), .ZN(net218284) );
  NAND2_X4 U6814 ( .A1(n5273), .A2(n5274), .ZN(n5525) );
  NAND2_X4 U6815 ( .A1(n5551), .A2(n5552), .ZN(n5624) );
  NAND2_X4 U6816 ( .A1(n5971), .A2(net215294), .ZN(net214730) );
  NAND2_X4 U6817 ( .A1(net216212), .A2(net216211), .ZN(net216020) );
  NAND2_X4 U6818 ( .A1(n5644), .A2(n5643), .ZN(n5508) );
  NAND2_X4 U6819 ( .A1(n7554), .A2(n7553), .ZN(n7374) );
  NAND2_X4 U6820 ( .A1(n3808), .A2(n5517), .ZN(net215809) );
  NAND2_X4 U6821 ( .A1(n5513), .A2(n5514), .ZN(n5772) );
  NAND2_X4 U6822 ( .A1(n3201), .A2(n6800), .ZN(n6884) );
  NAND2_X4 U6823 ( .A1(n7191), .A2(n7192), .ZN(net212652) );
  NAND2_X4 U6824 ( .A1(n7373), .A2(n7372), .ZN(n7553) );
  NAND2_X4 U6825 ( .A1(net213718), .A2(n6937), .ZN(net213594) );
  NAND2_X4 U6826 ( .A1(n6305), .A2(n3953), .ZN(n6383) );
  NAND2_X4 U6827 ( .A1(n3314), .A2(n5249), .ZN(n5480) );
  NAND2_X4 U6828 ( .A1(n5640), .A2(n5772), .ZN(n5515) );
  NAND2_X4 U6829 ( .A1(n5509), .A2(n3307), .ZN(n5803) );
  NAND2_X4 U6830 ( .A1(n4052), .A2(net218282), .ZN(net218097) );
  NAND3_X2 U6831 ( .A1(n5894), .A2(n5895), .A3(n5893), .ZN(n6149) );
  AOI21_X2 U6832 ( .B1(n3778), .B2(n5473), .A(n5345), .ZN(n5347) );
  INV_X2 U6833 ( .A(net216202), .ZN(net216198) );
  NAND2_X4 U6834 ( .A1(n4057), .A2(n4058), .ZN(net218267) );
  NAND2_X4 U6835 ( .A1(net212700), .A2(net212703), .ZN(n7204) );
  NAND2_X4 U6836 ( .A1(net213730), .A2(n6936), .ZN(net213581) );
  NAND2_X4 U6837 ( .A1(n7198), .A2(n7197), .ZN(net212954) );
  INV_X8 U6838 ( .A(n6609), .ZN(n6676) );
  NAND3_X2 U6839 ( .A1(a[1]), .A2(n5731), .A3(b[17]), .ZN(n5862) );
  NAND3_X1 U6840 ( .A1(n5305), .A2(n5304), .A3(n5618), .ZN(n5571) );
  NAND2_X1 U6841 ( .A1(n5304), .A2(n5618), .ZN(n5570) );
  NAND2_X1 U6842 ( .A1(n5078), .A2(n5080), .ZN(n5011) );
  OAI221_X1 U6843 ( .B1(net214479), .B2(net218600), .C1(n6625), .C2(n3991), 
        .A(net218610), .ZN(n6479) );
  NAND2_X4 U6844 ( .A1(n6832), .A2(n6833), .ZN(n6953) );
  NAND3_X2 U6845 ( .A1(a[0]), .A2(b[23]), .A3(n6625), .ZN(n6661) );
  NAND3_X1 U6846 ( .A1(n5909), .A2(n5910), .A3(n5908), .ZN(n5914) );
  AOI21_X2 U6847 ( .B1(n7236), .B2(n3926), .A(n7237), .ZN(n7199) );
  NOR2_X1 U6848 ( .A1(net218556), .A2(net219063), .ZN(n4298) );
  INV_X2 U6849 ( .A(n6787), .ZN(n6574) );
  NAND2_X4 U6850 ( .A1(n6787), .A2(n6786), .ZN(net214025) );
  NAND2_X4 U6851 ( .A1(n6507), .A2(n6506), .ZN(n6713) );
  NAND2_X4 U6852 ( .A1(net218658), .A2(a[0]), .ZN(net218655) );
  NAND2_X4 U6853 ( .A1(net218658), .A2(a[0]), .ZN(n3991) );
  NAND2_X4 U6854 ( .A1(net218658), .A2(a[0]), .ZN(n7888) );
  INV_X16 U6855 ( .A(net212094), .ZN(net212677) );
  NAND2_X4 U6856 ( .A1(net218548), .A2(net218544), .ZN(n7870) );
  INV_X32 U6857 ( .A(n3994), .ZN(n3995) );
  NAND2_X4 U6858 ( .A1(net218538), .A2(net218554), .ZN(n7871) );
  INV_X16 U6859 ( .A(n3995), .ZN(n7803) );
  INV_X16 U6860 ( .A(n7079), .ZN(n7039) );
  NAND2_X4 U6861 ( .A1(n7097), .A2(b[4]), .ZN(n4860) );
  INV_X32 U6862 ( .A(net218639), .ZN(net218640) );
  NAND2_X4 U6863 ( .A1(net217344), .A2(n4196), .ZN(net211994) );
  NAND2_X4 U6864 ( .A1(n7803), .A2(n4235), .ZN(n5330) );
  NAND2_X4 U6865 ( .A1(n7039), .A2(n4235), .ZN(n4942) );
  INV_X16 U6866 ( .A(n3993), .ZN(n7805) );
  NAND2_X4 U6867 ( .A1(n7805), .A2(n4235), .ZN(n5332) );
  NAND2_X4 U6868 ( .A1(n5446), .A2(n7039), .ZN(n6135) );
  INV_X16 U6869 ( .A(n6135), .ZN(n7050) );
  NAND2_X4 U6870 ( .A1(n4861), .A2(a[31]), .ZN(n7036) );
  INV_X16 U6871 ( .A(n3990), .ZN(n7389) );
  INV_X32 U6872 ( .A(net218628), .ZN(net218624) );
  INV_X32 U6873 ( .A(net218628), .ZN(net218626) );
  INV_X32 U6874 ( .A(net212283), .ZN(net218628) );
  INV_X32 U6875 ( .A(n3999), .ZN(n3997) );
  INV_X32 U6876 ( .A(n3999), .ZN(n3998) );
  INV_X32 U6877 ( .A(net218614), .ZN(net218606) );
  INV_X32 U6878 ( .A(net218614), .ZN(net218608) );
  INV_X32 U6879 ( .A(net218614), .ZN(net218610) );
  INV_X32 U6880 ( .A(net218604), .ZN(net218598) );
  INV_X32 U6881 ( .A(net218604), .ZN(net218600) );
  INV_X32 U6882 ( .A(b[1]), .ZN(net218566) );
  INV_X4 U6883 ( .A(op[0]), .ZN(net217346) );
  INV_X4 U6884 ( .A(op[2]), .ZN(net218371) );
  NAND4_X2 U6885 ( .A1(net218370), .A2(net218371), .A3(op[1]), .A4(op[0]), 
        .ZN(n4003) );
  NAND2_X2 U6886 ( .A1(n5193), .A2(b[9]), .ZN(n4167) );
  NAND2_X2 U6887 ( .A1(b[6]), .A2(a[2]), .ZN(n4141) );
  INV_X4 U6888 ( .A(n4141), .ZN(n4117) );
  OAI21_X4 U6889 ( .B1(net218362), .B2(net218352), .A(n4033), .ZN(n4120) );
  INV_X4 U6890 ( .A(n4017), .ZN(n4674) );
  NAND2_X2 U6891 ( .A1(n3343), .A2(n4674), .ZN(n4119) );
  XNOR2_X2 U6892 ( .A(n4067), .B(n4484), .ZN(n4009) );
  INV_X4 U6893 ( .A(n4009), .ZN(n4007) );
  XNOR2_X2 U6894 ( .A(n4005), .B(n4006), .ZN(n4025) );
  INV_X4 U6895 ( .A(n4028), .ZN(n4008) );
  NAND2_X2 U6896 ( .A1(a[3]), .A2(net218576), .ZN(net217654) );
  NAND2_X2 U6897 ( .A1(net218548), .A2(a[3]), .ZN(n4013) );
  INV_X4 U6898 ( .A(n4013), .ZN(n4014) );
  OAI211_X2 U6899 ( .C1(n4016), .C2(n3763), .A(n4015), .B(n4014), .ZN(
        net218217) );
  NAND3_X4 U6900 ( .A1(a[0]), .A2(a[1]), .A3(net218334), .ZN(n4026) );
  INV_X4 U6901 ( .A(n4248), .ZN(n4035) );
  XNOR2_X2 U6902 ( .A(n4031), .B(n4030), .ZN(net218273) );
  NAND2_X2 U6903 ( .A1(net218538), .A2(a[1]), .ZN(n4042) );
  INV_X4 U6904 ( .A(n4042), .ZN(n4040) );
  NOR3_X4 U6905 ( .A1(n4306), .A2(net218496), .A3(net218544), .ZN(n4058) );
  XNOR2_X2 U6906 ( .A(n4043), .B(n4042), .ZN(n4044) );
  XNOR2_X2 U6907 ( .A(n4044), .B(net220397), .ZN(n4057) );
  INV_X4 U6908 ( .A(n4045), .ZN(n4055) );
  NAND2_X2 U6909 ( .A1(net218550), .A2(net219055), .ZN(net218281) );
  INV_X4 U6910 ( .A(net218281), .ZN(net218282) );
  INV_X4 U6911 ( .A(n4050), .ZN(n4263) );
  NAND2_X2 U6912 ( .A1(n4263), .A2(n4049), .ZN(net218090) );
  NAND2_X2 U6913 ( .A1(net218090), .A2(n4068), .ZN(net218285) );
  XNOR2_X2 U6914 ( .A(net218284), .B(net218285), .ZN(n4053) );
  INV_X4 U6915 ( .A(net218266), .ZN(net218261) );
  NAND2_X2 U6916 ( .A1(b[4]), .A2(a[2]), .ZN(n4063) );
  OAI21_X4 U6917 ( .B1(net218262), .B2(net218263), .A(n4063), .ZN(n4092) );
  NOR2_X4 U6918 ( .A1(net218260), .A2(net218261), .ZN(n4056) );
  INV_X4 U6919 ( .A(net218251), .ZN(net218256) );
  XNOR2_X2 U6920 ( .A(n4056), .B(net218256), .ZN(n4079) );
  INV_X4 U6921 ( .A(n4079), .ZN(n4077) );
  NAND2_X2 U6922 ( .A1(b[4]), .A2(a[1]), .ZN(n4078) );
  XNOR2_X2 U6923 ( .A(n4059), .B(n4058), .ZN(n4328) );
  NAND3_X4 U6924 ( .A1(n4328), .A2(b[4]), .A3(a[0]), .ZN(n4087) );
  NAND2_X2 U6925 ( .A1(net218251), .A2(n4078), .ZN(n4060) );
  OAI21_X4 U6926 ( .B1(n4077), .B2(n4078), .A(n4062), .ZN(n4093) );
  INV_X4 U6927 ( .A(n4063), .ZN(n4064) );
  OAI21_X4 U6928 ( .B1(n4066), .B2(n4065), .A(net224032), .ZN(n4106) );
  INV_X4 U6929 ( .A(n4106), .ZN(n4075) );
  NAND2_X2 U6930 ( .A1(net218538), .A2(net219055), .ZN(net218210) );
  NAND2_X2 U6931 ( .A1(net218091), .A2(net218090), .ZN(net218232) );
  INV_X4 U6932 ( .A(net218232), .ZN(net218166) );
  INV_X4 U6933 ( .A(n4068), .ZN(n4069) );
  NOR3_X4 U6934 ( .A1(n4071), .A2(n4070), .A3(n4069), .ZN(n4122) );
  NAND2_X2 U6935 ( .A1(net218562), .A2(a[6]), .ZN(n4104) );
  XNOR2_X2 U6936 ( .A(n4104), .B(n4485), .ZN(net218165) );
  INV_X4 U6937 ( .A(n4072), .ZN(n4073) );
  INV_X4 U6938 ( .A(net218208), .ZN(net218207) );
  XNOR2_X2 U6939 ( .A(net218206), .B(net218207), .ZN(n4094) );
  NAND2_X2 U6940 ( .A1(a[3]), .A2(b[4]), .ZN(n4101) );
  INV_X4 U6941 ( .A(n4101), .ZN(n4095) );
  NAND2_X2 U6942 ( .A1(n4096), .A2(net218143), .ZN(n4074) );
  XNOR2_X2 U6943 ( .A(n4075), .B(n4074), .ZN(n4076) );
  NAND2_X2 U6944 ( .A1(b[5]), .A2(a[2]), .ZN(n4091) );
  NAND2_X2 U6945 ( .A1(n4077), .A2(n4078), .ZN(n4085) );
  INV_X4 U6946 ( .A(n4078), .ZN(n4080) );
  NAND2_X2 U6947 ( .A1(n4080), .A2(n4079), .ZN(n4086) );
  XNOR2_X2 U6948 ( .A(n4081), .B(n4087), .ZN(n4082) );
  NAND3_X4 U6949 ( .A1(b[5]), .A2(a[0]), .A3(n4380), .ZN(n4111) );
  INV_X4 U6950 ( .A(n4111), .ZN(n4084) );
  NAND2_X2 U6951 ( .A1(b[5]), .A2(a[1]), .ZN(n4107) );
  NAND2_X2 U6952 ( .A1(n4108), .A2(n4107), .ZN(n4083) );
  INV_X4 U6953 ( .A(n4107), .ZN(n4090) );
  XNOR2_X2 U6954 ( .A(n4109), .B(n4108), .ZN(n4089) );
  INV_X4 U6955 ( .A(net218041), .ZN(net218178) );
  INV_X4 U6956 ( .A(n4091), .ZN(n4100) );
  XNOR2_X2 U6957 ( .A(n4098), .B(n4097), .ZN(n4099) );
  NAND3_X4 U6958 ( .A1(net218143), .A2(net224032), .A3(net218116), .ZN(
        net217240) );
  INV_X4 U6959 ( .A(n4104), .ZN(n4105) );
  NAND2_X2 U6960 ( .A1(n4359), .A2(n4105), .ZN(net218089) );
  NAND2_X2 U6961 ( .A1(net218548), .A2(a[6]), .ZN(net218157) );
  XNOR2_X2 U6962 ( .A(net218149), .B(net217244), .ZN(net218144) );
  NAND2_X2 U6963 ( .A1(a[3]), .A2(b[5]), .ZN(net218137) );
  XNOR2_X2 U6964 ( .A(net218132), .B(net218133), .ZN(n4140) );
  XNOR2_X2 U6965 ( .A(n4108), .B(n4107), .ZN(n4110) );
  XNOR2_X2 U6966 ( .A(n4110), .B(n4109), .ZN(n4112) );
  XNOR2_X2 U6967 ( .A(n4112), .B(n4111), .ZN(n4410) );
  NAND2_X2 U6968 ( .A1(b[6]), .A2(a[1]), .ZN(n4145) );
  INV_X4 U6969 ( .A(n4145), .ZN(n4135) );
  XNOR2_X2 U6970 ( .A(net218124), .B(net218041), .ZN(n4114) );
  OAI21_X4 U6971 ( .B1(n4115), .B2(n4114), .A(n4113), .ZN(n4116) );
  OAI21_X4 U6972 ( .B1(n4117), .B2(n3935), .A(n4116), .ZN(n4793) );
  INV_X4 U6973 ( .A(net217244), .ZN(net217732) );
  NAND2_X2 U6974 ( .A1(net218548), .A2(a[7]), .ZN(n4123) );
  INV_X4 U6975 ( .A(net217141), .ZN(net218084) );
  INV_X4 U6976 ( .A(net218076), .ZN(net218075) );
  NAND3_X4 U6977 ( .A1(net218075), .A2(a[7]), .A3(net218546), .ZN(n4798) );
  XNOR2_X2 U6978 ( .A(n4125), .B(n4124), .ZN(net217284) );
  NAND2_X2 U6979 ( .A1(net218538), .A2(a[6]), .ZN(net217285) );
  NAND2_X2 U6980 ( .A1(a[3]), .A2(b[6]), .ZN(n4126) );
  INV_X4 U6981 ( .A(n4126), .ZN(n4128) );
  XNOR2_X2 U6982 ( .A(n4731), .B(n4129), .ZN(n4132) );
  INV_X4 U6983 ( .A(n4132), .ZN(n4130) );
  NAND2_X2 U6984 ( .A1(b[7]), .A2(a[2]), .ZN(n4131) );
  INV_X4 U6985 ( .A(n4131), .ZN(n4133) );
  NAND2_X2 U6986 ( .A1(n4133), .A2(n4132), .ZN(n4741) );
  NAND2_X2 U6987 ( .A1(n4735), .A2(n4741), .ZN(n4157) );
  XNOR2_X2 U6988 ( .A(net218040), .B(net218041), .ZN(n4134) );
  NAND2_X2 U6989 ( .A1(n4146), .A2(n4145), .ZN(n4138) );
  INV_X4 U6990 ( .A(n4152), .ZN(n4136) );
  AOI21_X4 U6991 ( .B1(n4138), .B2(n4137), .A(n4136), .ZN(n4139) );
  XNOR2_X2 U6992 ( .A(n4139), .B(n3316), .ZN(n4144) );
  INV_X4 U6993 ( .A(n4140), .ZN(n4142) );
  XNOR2_X2 U6994 ( .A(n4144), .B(n4143), .ZN(n4739) );
  INV_X4 U6995 ( .A(n4739), .ZN(n4163) );
  NAND2_X2 U6996 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  XNOR2_X2 U6997 ( .A(n4148), .B(n4151), .ZN(n4149) );
  INV_X4 U6998 ( .A(n4149), .ZN(n4444) );
  NAND3_X4 U6999 ( .A1(b[7]), .A2(a[0]), .A3(n4444), .ZN(n4737) );
  XNOR2_X2 U7000 ( .A(n4154), .B(n4153), .ZN(n4155) );
  XNOR2_X2 U7001 ( .A(n4157), .B(n4156), .ZN(n4160) );
  NAND2_X2 U7002 ( .A1(b[8]), .A2(a[1]), .ZN(n4159) );
  INV_X4 U7003 ( .A(n4159), .ZN(n4161) );
  NAND2_X2 U7004 ( .A1(n4161), .A2(n4160), .ZN(n4825) );
  INV_X4 U7005 ( .A(n4737), .ZN(n4162) );
  XNOR2_X2 U7006 ( .A(n4163), .B(n4162), .ZN(n4477) );
  XNOR2_X2 U7007 ( .A(n4164), .B(n4824), .ZN(n4165) );
  INV_X4 U7008 ( .A(n4165), .ZN(n4754) );
  MUX2_X2 U7009 ( .A(n4167), .B(n4166), .S(n4754), .Z(n4202) );
  INV_X4 U7010 ( .A(op[2]), .ZN(net217946) );
  XNOR2_X2 U7011 ( .A(n4002), .B(b[7]), .ZN(n4175) );
  XNOR2_X2 U7012 ( .A(n4175), .B(net218442), .ZN(n4456) );
  XNOR2_X2 U7013 ( .A(sel), .B(b[5]), .ZN(n4174) );
  XNOR2_X2 U7014 ( .A(n4174), .B(net218456), .ZN(n4389) );
  XNOR2_X2 U7015 ( .A(sel), .B(net218534), .ZN(n4173) );
  XNOR2_X2 U7016 ( .A(sel), .B(net218558), .ZN(n4172) );
  XNOR2_X2 U7017 ( .A(n4172), .B(net218484), .ZN(n4256) );
  XNOR2_X2 U7018 ( .A(sel), .B(net218574), .ZN(n4168) );
  INV_X4 U7019 ( .A(n4168), .ZN(n4171) );
  XNOR2_X2 U7020 ( .A(n4168), .B(net218496), .ZN(n4695) );
  INV_X4 U7021 ( .A(n4695), .ZN(n4169) );
  NAND2_X2 U7022 ( .A1(n4000), .A2(n4169), .ZN(n4697) );
  INV_X4 U7023 ( .A(n4697), .ZN(n4170) );
  AOI21_X4 U7024 ( .B1(a[0]), .B2(n4171), .A(n4170), .ZN(n4257) );
  OAI22_X2 U7025 ( .A1(n4172), .A2(net218486), .B1(n4256), .B2(n4257), .ZN(
        n4203) );
  XNOR2_X2 U7026 ( .A(n4000), .B(net218546), .ZN(net217995) );
  INV_X4 U7027 ( .A(net217933), .ZN(net217993) );
  INV_X4 U7028 ( .A(net217995), .ZN(net217994) );
  AOI22_X2 U7029 ( .A1(n4203), .A2(net217993), .B1(a[2]), .B2(net217994), .ZN(
        n4295) );
  XNOR2_X2 U7030 ( .A(sel), .B(b[4]), .ZN(net217990) );
  INV_X4 U7031 ( .A(net217761), .ZN(net217988) );
  INV_X4 U7032 ( .A(net217990), .ZN(net217989) );
  AOI22_X2 U7033 ( .A1(n4332), .A2(net217988), .B1(net219055), .B2(net217989), 
        .ZN(n4390) );
  OAI22_X2 U7034 ( .A1(n4174), .A2(net218456), .B1(n4389), .B2(n4390), .ZN(
        n4424) );
  XNOR2_X2 U7035 ( .A(n4000), .B(b[6]), .ZN(net217984) );
  INV_X4 U7036 ( .A(n3354), .ZN(net217982) );
  INV_X4 U7037 ( .A(net217984), .ZN(net217983) );
  AOI22_X2 U7038 ( .A1(n4424), .A2(net217982), .B1(a[6]), .B2(net217983), .ZN(
        n4457) );
  OAI22_X2 U7039 ( .A1(n4175), .A2(net218442), .B1(n4456), .B2(n4457), .ZN(
        n4481) );
  XNOR2_X2 U7040 ( .A(sel), .B(b[8]), .ZN(net217979) );
  INV_X4 U7041 ( .A(net217584), .ZN(net217977) );
  INV_X4 U7042 ( .A(net217979), .ZN(net217978) );
  AOI22_X2 U7043 ( .A1(n4481), .A2(net217977), .B1(a[8]), .B2(net217978), .ZN(
        n4760) );
  XNOR2_X2 U7044 ( .A(n4000), .B(b[9]), .ZN(n4761) );
  XNOR2_X2 U7045 ( .A(n4761), .B(net218428), .ZN(n4759) );
  INV_X4 U7046 ( .A(n4759), .ZN(n4176) );
  XNOR2_X2 U7047 ( .A(n4760), .B(n4176), .ZN(n4189) );
  NAND2_X2 U7048 ( .A1(net218578), .A2(net218566), .ZN(n4177) );
  INV_X4 U7049 ( .A(n4177), .ZN(n7855) );
  NAND2_X2 U7050 ( .A1(n3997), .A2(a[5]), .ZN(net217860) );
  INV_X4 U7051 ( .A(net217860), .ZN(net217973) );
  INV_X4 U7052 ( .A(net217759), .ZN(net212283) );
  NAND2_X2 U7053 ( .A1(net218626), .A2(a[3]), .ZN(n4264) );
  INV_X4 U7054 ( .A(n4264), .ZN(n4178) );
  NOR2_X4 U7055 ( .A1(net217973), .A2(n4178), .ZN(n4179) );
  NAND2_X2 U7056 ( .A1(n4179), .A2(net217972), .ZN(n5595) );
  INV_X4 U7057 ( .A(n5595), .ZN(n6102) );
  NAND2_X2 U7058 ( .A1(n3997), .A2(a[1]), .ZN(n4267) );
  NAND2_X2 U7059 ( .A1(n7803), .A2(n6100), .ZN(n4181) );
  NAND2_X2 U7060 ( .A1(net218554), .A2(net218544), .ZN(n7079) );
  NAND2_X2 U7061 ( .A1(n4263), .A2(net218556), .ZN(n4297) );
  NAND2_X2 U7062 ( .A1(net218626), .A2(a[7]), .ZN(net217859) );
  NAND2_X2 U7063 ( .A1(n3997), .A2(a[9]), .ZN(net217942) );
  NAND4_X2 U7064 ( .A1(net217816), .A2(n4297), .A3(net217859), .A4(net217942), 
        .ZN(n6123) );
  NAND2_X2 U7065 ( .A1(n7039), .A2(n6123), .ZN(n4180) );
  OAI211_X2 U7066 ( .C1(n6102), .C2(n3993), .A(n4181), .B(n4180), .ZN(n4182)
         );
  INV_X4 U7067 ( .A(n4182), .ZN(n6861) );
  NOR2_X4 U7068 ( .A1(op[0]), .A2(op[1]), .ZN(n4183) );
  INV_X4 U7069 ( .A(net217966), .ZN(net217950) );
  NAND2_X2 U7070 ( .A1(n4183), .A2(net217950), .ZN(n7878) );
  INV_X4 U7071 ( .A(n7878), .ZN(n7821) );
  NAND2_X2 U7072 ( .A1(n7821), .A2(net218530), .ZN(n5323) );
  NAND2_X2 U7073 ( .A1(n3997), .A2(a[29]), .ZN(n7215) );
  INV_X4 U7074 ( .A(n7438), .ZN(n7436) );
  NAND2_X2 U7075 ( .A1(n7436), .A2(net218566), .ZN(n7865) );
  NAND2_X2 U7076 ( .A1(n7215), .A2(n7865), .ZN(n4184) );
  INV_X4 U7077 ( .A(n4184), .ZN(n4191) );
  NAND2_X2 U7078 ( .A1(a[31]), .A2(net218558), .ZN(n4185) );
  NAND2_X2 U7079 ( .A1(n4191), .A2(n4185), .ZN(n5054) );
  INV_X4 U7080 ( .A(n5054), .ZN(n7381) );
  NAND2_X2 U7081 ( .A1(a[31]), .A2(net218538), .ZN(n6636) );
  NAND2_X2 U7082 ( .A1(a[26]), .A2(net218574), .ZN(net213830) );
  NAND2_X2 U7083 ( .A1(net217782), .A2(net218566), .ZN(net213330) );
  INV_X4 U7084 ( .A(n7217), .ZN(n4186) );
  NAND2_X2 U7085 ( .A1(n4186), .A2(net218556), .ZN(n7864) );
  NAND2_X2 U7086 ( .A1(net218626), .A2(a[27]), .ZN(n7216) );
  NAND2_X2 U7087 ( .A1(n3997), .A2(a[25]), .ZN(net213927) );
  NAND4_X2 U7088 ( .A1(net213330), .A2(n7864), .A3(n7216), .A4(net213927), 
        .ZN(n4383) );
  NAND2_X2 U7089 ( .A1(n7039), .A2(n4383), .ZN(n4192) );
  OAI211_X2 U7090 ( .C1(n7381), .C2(n3993), .A(n6636), .B(n4192), .ZN(n6855)
         );
  INV_X4 U7091 ( .A(n6855), .ZN(n4187) );
  NAND2_X2 U7092 ( .A1(net217960), .A2(net217950), .ZN(n4673) );
  INV_X4 U7093 ( .A(n4673), .ZN(n7858) );
  NAND2_X2 U7094 ( .A1(n7858), .A2(b[4]), .ZN(n4768) );
  OAI22_X2 U7095 ( .A1(n6861), .A2(n5323), .B1(n4187), .B2(n4768), .ZN(n4188)
         );
  AOI21_X2 U7096 ( .B1(n4189), .B2(n3990), .A(n4188), .ZN(n4201) );
  NAND2_X2 U7097 ( .A1(net218626), .A2(a[31]), .ZN(n4190) );
  NAND2_X2 U7098 ( .A1(n4191), .A2(n4190), .ZN(n7380) );
  INV_X4 U7099 ( .A(n7380), .ZN(n4193) );
  INV_X4 U7100 ( .A(n4194), .ZN(n6845) );
  NOR2_X4 U7101 ( .A1(op[1]), .A2(net217346), .ZN(n4195) );
  NAND2_X2 U7102 ( .A1(net217950), .A2(n4195), .ZN(n4672) );
  INV_X4 U7103 ( .A(n4672), .ZN(n7097) );
  INV_X4 U7104 ( .A(net217948), .ZN(net217344) );
  NOR2_X4 U7105 ( .A1(op[0]), .A2(op[2]), .ZN(n4196) );
  INV_X4 U7106 ( .A(net217944), .ZN(net217943) );
  NOR2_X4 U7107 ( .A1(b[9]), .A2(a[9]), .ZN(n4508) );
  NAND2_X2 U7108 ( .A1(a[18]), .A2(net218576), .ZN(net215853) );
  NAND2_X2 U7109 ( .A1(net217807), .A2(net218566), .ZN(net215491) );
  NAND2_X2 U7110 ( .A1(a[20]), .A2(net218574), .ZN(net215421) );
  NAND2_X2 U7111 ( .A1(net218626), .A2(a[19]), .ZN(n6114) );
  NAND2_X2 U7112 ( .A1(n3997), .A2(a[17]), .ZN(n5596) );
  NAND4_X2 U7113 ( .A1(net215491), .A2(net214487), .A3(n6114), .A4(n5596), 
        .ZN(n4279) );
  INV_X4 U7114 ( .A(n4279), .ZN(n5058) );
  NAND2_X2 U7115 ( .A1(n7097), .A2(net218530), .ZN(n7035) );
  NAND2_X2 U7116 ( .A1(n7858), .A2(net218530), .ZN(n6637) );
  NAND2_X2 U7117 ( .A1(n7035), .A2(n6637), .ZN(n4235) );
  OAI222_X2 U7118 ( .A1(n6845), .A2(n4860), .B1(net217943), .B2(n4508), .C1(
        n5058), .C2(n5330), .ZN(n4199) );
  NAND2_X2 U7119 ( .A1(net218626), .A2(a[11]), .ZN(net216710) );
  NAND2_X2 U7120 ( .A1(net218576), .A2(a[12]), .ZN(net216965) );
  NAND2_X2 U7121 ( .A1(net217818), .A2(net218558), .ZN(net216328) );
  INV_X4 U7122 ( .A(net217271), .ZN(net217817) );
  NAND2_X2 U7123 ( .A1(net217817), .A2(net218566), .ZN(net217027) );
  NAND2_X2 U7124 ( .A1(a[22]), .A2(net218574), .ZN(net214926) );
  NAND2_X2 U7125 ( .A1(net217780), .A2(net218566), .ZN(net214486) );
  NAND2_X2 U7126 ( .A1(a[24]), .A2(net218574), .ZN(net214391) );
  NAND2_X2 U7127 ( .A1(net217783), .A2(net218558), .ZN(net213331) );
  NAND2_X2 U7128 ( .A1(net218626), .A2(a[23]), .ZN(net213926) );
  NAND2_X2 U7129 ( .A1(n3997), .A2(a[21]), .ZN(net215024) );
  INV_X4 U7130 ( .A(net217838), .ZN(net216692) );
  NAND2_X2 U7131 ( .A1(net218538), .A2(net218550), .ZN(n7869) );
  NAND2_X2 U7132 ( .A1(n3997), .A2(a[13]), .ZN(net216711) );
  NAND2_X2 U7133 ( .A1(net218576), .A2(a[16]), .ZN(net216256) );
  NAND2_X2 U7134 ( .A1(net217806), .A2(net218558), .ZN(net215492) );
  NAND2_X2 U7135 ( .A1(net218626), .A2(a[15]), .ZN(net215920) );
  NAND2_X2 U7136 ( .A1(a[14]), .A2(net218576), .ZN(net216627) );
  INV_X4 U7137 ( .A(net216627), .ZN(net217819) );
  NAND2_X2 U7138 ( .A1(net217819), .A2(net218566), .ZN(net216327) );
  INV_X4 U7139 ( .A(net216704), .ZN(net217849) );
  OAI22_X2 U7140 ( .A1(net216692), .A2(n3996), .B1(net217849), .B2(n5332), 
        .ZN(n4197) );
  NOR3_X4 U7141 ( .A1(n4199), .A2(n4198), .A3(n4197), .ZN(n4200) );
  NAND4_X2 U7142 ( .A1(n4202), .A2(n3397), .A3(n4201), .A4(n4200), .ZN(
        result[9]) );
  XNOR2_X2 U7143 ( .A(n4203), .B(net217933), .ZN(n4209) );
  MUX2_X2 U7144 ( .A(net217654), .B(n3909), .S(net218560), .Z(n4204) );
  INV_X4 U7145 ( .A(n4204), .ZN(n4206) );
  NAND2_X2 U7146 ( .A1(n3997), .A2(a[2]), .ZN(n4242) );
  NAND2_X2 U7147 ( .A1(n4418), .A2(n4242), .ZN(n4205) );
  AOI21_X2 U7148 ( .B1(n4209), .B2(n3990), .A(n4208), .ZN(n4255) );
  INV_X4 U7149 ( .A(n4860), .ZN(n5051) );
  NAND2_X2 U7150 ( .A1(net218626), .A2(a[24]), .ZN(n4210) );
  INV_X4 U7151 ( .A(n4210), .ZN(n6992) );
  NOR2_X4 U7152 ( .A1(n6992), .A2(n3368), .ZN(n4212) );
  MUX2_X2 U7153 ( .A(net213634), .B(net213311), .S(net218558), .Z(n4211) );
  NAND2_X2 U7154 ( .A1(n4212), .A2(n4211), .ZN(n4778) );
  NAND2_X2 U7155 ( .A1(n7805), .A2(n4778), .ZN(n4221) );
  NAND2_X2 U7156 ( .A1(net218626), .A2(a[20]), .ZN(n4213) );
  INV_X4 U7157 ( .A(n4213), .ZN(n6132) );
  NOR2_X4 U7158 ( .A1(n6132), .A2(n3367), .ZN(n4215) );
  NAND2_X2 U7159 ( .A1(a[19]), .A2(net218574), .ZN(net215001) );
  MUX2_X2 U7160 ( .A(net215001), .B(net214224), .S(net218556), .Z(n4214) );
  NAND2_X2 U7161 ( .A1(n4215), .A2(n4214), .ZN(n4774) );
  NAND2_X2 U7162 ( .A1(n7039), .A2(n4774), .ZN(n4220) );
  NAND2_X2 U7163 ( .A1(net218626), .A2(a[28]), .ZN(n4216) );
  INV_X4 U7164 ( .A(n4216), .ZN(n7815) );
  NOR2_X4 U7165 ( .A1(n3371), .A2(n7815), .ZN(n4218) );
  MUX2_X2 U7166 ( .A(n7816), .B(n7817), .S(net218558), .Z(n4217) );
  NAND2_X2 U7167 ( .A1(n4218), .A2(n4217), .ZN(n5178) );
  NAND2_X2 U7168 ( .A1(n7803), .A2(n5178), .ZN(n4219) );
  INV_X4 U7169 ( .A(n4241), .ZN(n4224) );
  NAND2_X2 U7170 ( .A1(n3997), .A2(a[30]), .ZN(n7813) );
  INV_X4 U7171 ( .A(n7668), .ZN(n4222) );
  NAND2_X2 U7172 ( .A1(n4222), .A2(net218566), .ZN(n7669) );
  NAND2_X2 U7173 ( .A1(n7813), .A2(n7669), .ZN(n7831) );
  NAND2_X2 U7174 ( .A1(n7807), .A2(n7831), .ZN(n4223) );
  NAND2_X2 U7175 ( .A1(n4224), .A2(n4223), .ZN(n5745) );
  NAND2_X2 U7176 ( .A1(n5051), .A2(n5745), .ZN(n4254) );
  NAND2_X2 U7177 ( .A1(net218626), .A2(a[16]), .ZN(n4225) );
  INV_X4 U7178 ( .A(n4225), .ZN(n5746) );
  NOR2_X4 U7179 ( .A1(n5746), .A2(n3366), .ZN(n4227) );
  NAND2_X2 U7180 ( .A1(net218574), .A2(a[15]), .ZN(net215701) );
  MUX2_X2 U7181 ( .A(net215701), .B(net215245), .S(net218558), .Z(n4226) );
  NAND2_X2 U7182 ( .A1(n4227), .A2(n4226), .ZN(n5167) );
  INV_X4 U7183 ( .A(n5167), .ZN(n4779) );
  NOR2_X4 U7184 ( .A1(net218546), .A2(a[2]), .ZN(n4244) );
  NAND2_X2 U7185 ( .A1(net218624), .A2(a[12]), .ZN(n4228) );
  INV_X4 U7186 ( .A(n4228), .ZN(n5162) );
  NAND2_X2 U7187 ( .A1(n3997), .A2(a[10]), .ZN(n4764) );
  INV_X4 U7188 ( .A(n4764), .ZN(n4229) );
  NOR2_X4 U7189 ( .A1(n5162), .A2(n4229), .ZN(n4231) );
  MUX2_X2 U7190 ( .A(net216517), .B(net216117), .S(net218556), .Z(n4230) );
  NAND2_X2 U7191 ( .A1(n4231), .A2(n4230), .ZN(n4427) );
  NAND2_X2 U7192 ( .A1(n7803), .A2(n4427), .ZN(n4237) );
  INV_X4 U7193 ( .A(net217182), .ZN(net217897) );
  NAND2_X2 U7194 ( .A1(n3997), .A2(a[6]), .ZN(n4232) );
  INV_X4 U7195 ( .A(n4232), .ZN(n4420) );
  NOR2_X4 U7196 ( .A1(net217897), .A2(n4420), .ZN(n4234) );
  MUX2_X2 U7197 ( .A(n4485), .B(net216885), .S(net218558), .Z(n4233) );
  NAND2_X2 U7198 ( .A1(n4234), .A2(n4233), .ZN(n4432) );
  NAND2_X2 U7199 ( .A1(n7805), .A2(n4432), .ZN(n4236) );
  INV_X4 U7200 ( .A(n4235), .ZN(n6653) );
  NOR3_X4 U7201 ( .A1(n4240), .A2(n4239), .A3(n4238), .ZN(n4253) );
  INV_X4 U7202 ( .A(a[31]), .ZN(net217557) );
  OAI21_X4 U7203 ( .B1(n3997), .B2(net217557), .A(n7813), .ZN(n7829) );
  AOI21_X4 U7204 ( .B1(n7807), .B2(n7829), .A(n4241), .ZN(n5750) );
  INV_X4 U7205 ( .A(n5323), .ZN(n5446) );
  NAND2_X2 U7206 ( .A1(net218624), .A2(a[0]), .ZN(n4243) );
  NAND2_X2 U7207 ( .A1(net218576), .A2(a[1]), .ZN(n4349) );
  INV_X4 U7208 ( .A(n4349), .ZN(n4274) );
  NAND2_X2 U7209 ( .A1(n4274), .A2(net218566), .ZN(n4677) );
  NAND3_X2 U7210 ( .A1(n4243), .A2(n4242), .A3(n4677), .ZN(n6272) );
  NAND2_X2 U7211 ( .A1(n7050), .A2(n6272), .ZN(n4247) );
  INV_X4 U7212 ( .A(n4244), .ZN(n4245) );
  NAND2_X2 U7213 ( .A1(n4245), .A2(n4248), .ZN(n4582) );
  INV_X4 U7214 ( .A(n4582), .ZN(n4600) );
  NAND2_X2 U7215 ( .A1(n4600), .A2(net218639), .ZN(n4246) );
  OAI211_X2 U7216 ( .C1(n5750), .C2(n4768), .A(n4247), .B(n4246), .ZN(n4251)
         );
  NAND2_X2 U7217 ( .A1(net218658), .A2(net218554), .ZN(n4249) );
  NAND2_X2 U7218 ( .A1(n4249), .A2(net212094), .ZN(net217878) );
  NOR3_X2 U7219 ( .A1(n4251), .A2(n4250), .A3(net217876), .ZN(n4252) );
  NAND4_X2 U7220 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(
        result[2]) );
  INV_X4 U7221 ( .A(n4256), .ZN(n4258) );
  XNOR2_X2 U7222 ( .A(n4258), .B(n4257), .ZN(n4261) );
  NAND2_X2 U7223 ( .A1(n7050), .A2(n6100), .ZN(n4259) );
  INV_X4 U7224 ( .A(n4259), .ZN(n4260) );
  AOI21_X2 U7225 ( .B1(n4261), .B2(n3990), .A(n4260), .ZN(n4293) );
  INV_X4 U7226 ( .A(net217433), .ZN(net217545) );
  NAND2_X2 U7227 ( .A1(net217545), .A2(net218639), .ZN(n4292) );
  NAND2_X2 U7228 ( .A1(n4263), .A2(net218566), .ZN(net217621) );
  INV_X4 U7229 ( .A(net217858), .ZN(net217677) );
  NAND2_X2 U7230 ( .A1(n4265), .A2(n4264), .ZN(n4269) );
  NAND2_X2 U7231 ( .A1(n4267), .A2(n4449), .ZN(n4268) );
  OAI21_X4 U7232 ( .B1(net217677), .B2(n3993), .A(n4270), .ZN(n4273) );
  NOR2_X4 U7233 ( .A1(n3360), .A2(n3995), .ZN(n4272) );
  NOR2_X4 U7234 ( .A1(net217849), .A2(n7869), .ZN(n4271) );
  NOR3_X4 U7235 ( .A1(n4273), .A2(n4272), .A3(n4271), .ZN(n4278) );
  OAI211_X2 U7236 ( .C1(n4274), .C2(n3991), .A(net211950), .B(n3411), .ZN(
        n4276) );
  AOI21_X2 U7237 ( .B1(net218556), .B2(n4276), .A(n4275), .ZN(n4277) );
  OAI21_X4 U7238 ( .B1(n6653), .B2(n4278), .A(n4277), .ZN(n4289) );
  NAND2_X2 U7239 ( .A1(n7803), .A2(n4383), .ZN(n4282) );
  NAND2_X2 U7240 ( .A1(n7805), .A2(net217838), .ZN(n4281) );
  NAND2_X2 U7241 ( .A1(n7039), .A2(n4279), .ZN(n4280) );
  NAND3_X2 U7242 ( .A1(n4282), .A2(n4281), .A3(n4280), .ZN(n4286) );
  INV_X4 U7243 ( .A(n4286), .ZN(n4284) );
  NAND2_X2 U7244 ( .A1(n7807), .A2(n7380), .ZN(n4283) );
  NAND2_X2 U7245 ( .A1(n4284), .A2(n4283), .ZN(n5602) );
  INV_X4 U7246 ( .A(n5602), .ZN(n4285) );
  NOR2_X4 U7247 ( .A1(n4285), .A2(n4860), .ZN(n4288) );
  AOI21_X4 U7248 ( .B1(n7807), .B2(n5054), .A(n4286), .ZN(n5607) );
  NOR2_X4 U7249 ( .A1(n5607), .A2(n4768), .ZN(n4287) );
  NOR3_X4 U7250 ( .A1(n4289), .A2(n4288), .A3(n4287), .ZN(n4290) );
  NAND4_X2 U7251 ( .A1(n4293), .A2(n4292), .A3(n4291), .A4(n4290), .ZN(
        result[1]) );
  INV_X4 U7252 ( .A(n4294), .ZN(n4296) );
  XNOR2_X2 U7253 ( .A(n4296), .B(n4295), .ZN(n4304) );
  NAND2_X2 U7254 ( .A1(net218624), .A2(a[13]), .ZN(net216330) );
  NAND2_X2 U7255 ( .A1(net217819), .A2(net218558), .ZN(net215919) );
  NAND2_X2 U7256 ( .A1(net217818), .A2(net218566), .ZN(n5045) );
  NAND2_X2 U7257 ( .A1(n3997), .A2(a[11]), .ZN(net217030) );
  NAND4_X2 U7258 ( .A1(net216330), .A2(net215919), .A3(n5045), .A4(net217030), 
        .ZN(n4856) );
  INV_X4 U7259 ( .A(n4856), .ZN(n4460) );
  NAND2_X2 U7260 ( .A1(net218624), .A2(a[9]), .ZN(net217029) );
  NAND2_X2 U7261 ( .A1(n3998), .A2(a[7]), .ZN(n4447) );
  NOR2_X4 U7262 ( .A1(net218534), .A2(a[3]), .ZN(net217796) );
  OAI221_X2 U7263 ( .B1(n4460), .B2(n5330), .C1(n3333), .C2(n5332), .A(n3408), 
        .ZN(n4303) );
  NAND2_X2 U7264 ( .A1(net218624), .A2(a[5]), .ZN(n4448) );
  NAND2_X2 U7265 ( .A1(n3998), .A2(a[3]), .ZN(n4310) );
  NAND2_X2 U7266 ( .A1(n4448), .A2(n4310), .ZN(n4300) );
  INV_X4 U7267 ( .A(n4297), .ZN(n4299) );
  NAND2_X2 U7268 ( .A1(n3998), .A2(a[15]), .ZN(net216329) );
  NAND2_X2 U7269 ( .A1(net217807), .A2(net218558), .ZN(net215023) );
  NAND2_X2 U7270 ( .A1(net217806), .A2(net218566), .ZN(n5597) );
  NAND2_X2 U7271 ( .A1(net218624), .A2(a[17]), .ZN(net215494) );
  NAND4_X2 U7272 ( .A1(net216329), .A2(net215023), .A3(n5597), .A4(net215494), 
        .ZN(n5320) );
  INV_X4 U7273 ( .A(n5320), .ZN(n4867) );
  OAI22_X2 U7274 ( .A1(n4301), .A2(n4942), .B1(n4867), .B2(n3996), .ZN(n4302)
         );
  AOI211_X2 U7275 ( .C1(n4304), .C2(n3990), .A(n4303), .B(n4302), .ZN(n4326)
         );
  NAND2_X2 U7276 ( .A1(net218658), .A2(net218544), .ZN(n4305) );
  NAND2_X2 U7277 ( .A1(n4305), .A2(net212094), .ZN(n4308) );
  INV_X4 U7278 ( .A(n4306), .ZN(n4307) );
  MUX2_X2 U7279 ( .A(n4309), .B(n4308), .S(n4307), .Z(n4324) );
  INV_X4 U7280 ( .A(net217796), .ZN(net217795) );
  INV_X4 U7281 ( .A(n4310), .ZN(n4312) );
  NOR2_X4 U7282 ( .A1(n4312), .A2(n4311), .ZN(n4314) );
  MUX2_X2 U7283 ( .A(n3881), .B(n4700), .S(net218556), .Z(n4313) );
  NAND2_X2 U7284 ( .A1(n4314), .A2(n4313), .ZN(n5315) );
  INV_X4 U7285 ( .A(n5315), .ZN(n6453) );
  NAND2_X2 U7286 ( .A1(n3998), .A2(a[27]), .ZN(net213332) );
  INV_X4 U7287 ( .A(net213332), .ZN(net217786) );
  NAND2_X2 U7288 ( .A1(net218624), .A2(a[29]), .ZN(n7862) );
  INV_X4 U7289 ( .A(n7862), .ZN(n4315) );
  NOR2_X4 U7290 ( .A1(net217786), .A2(n4315), .ZN(n4317) );
  MUX2_X2 U7291 ( .A(n7217), .B(n7438), .S(net218560), .Z(n4316) );
  NAND2_X2 U7292 ( .A1(n4317), .A2(n4316), .ZN(n4865) );
  INV_X4 U7293 ( .A(n4865), .ZN(n7041) );
  NAND2_X2 U7294 ( .A1(n3998), .A2(a[31]), .ZN(n7863) );
  MUX2_X2 U7295 ( .A(n7041), .B(n7863), .S(net218546), .Z(n7038) );
  NAND2_X2 U7296 ( .A1(net217783), .A2(net218566), .ZN(net213924) );
  NAND2_X2 U7297 ( .A1(net217782), .A2(net218556), .ZN(n6921) );
  NAND2_X2 U7298 ( .A1(n3998), .A2(a[23]), .ZN(n6470) );
  NAND2_X2 U7299 ( .A1(net218624), .A2(a[25]), .ZN(net213333) );
  NAND4_X2 U7300 ( .A1(net213924), .A2(n6921), .A3(n6470), .A4(net213333), 
        .ZN(n4450) );
  INV_X4 U7301 ( .A(n4450), .ZN(n5331) );
  NAND2_X2 U7302 ( .A1(net217781), .A2(net218566), .ZN(net215022) );
  NAND2_X2 U7303 ( .A1(net217780), .A2(net218556), .ZN(net213925) );
  NAND2_X2 U7304 ( .A1(n3998), .A2(a[19]), .ZN(net215493) );
  NAND2_X2 U7305 ( .A1(net218624), .A2(a[21]), .ZN(net214489) );
  INV_X4 U7306 ( .A(net217779), .ZN(net216306) );
  OAI22_X2 U7307 ( .A1(n5331), .A2(n3993), .B1(net216306), .B2(n7079), .ZN(
        n4318) );
  INV_X4 U7308 ( .A(n4318), .ZN(n4320) );
  INV_X4 U7309 ( .A(n4319), .ZN(n5880) );
  INV_X4 U7310 ( .A(n4768), .ZN(n4861) );
  NAND2_X2 U7311 ( .A1(n7807), .A2(a[31]), .ZN(n4416) );
  OAI211_X2 U7312 ( .C1(n7041), .C2(n3995), .A(n4416), .B(n4320), .ZN(n5877)
         );
  NAND2_X2 U7313 ( .A1(n4861), .A2(n5877), .ZN(n4321) );
  NOR4_X2 U7314 ( .A1(n4324), .A2(net217771), .A3(n4323), .A4(n4322), .ZN(
        n4325) );
  NAND2_X2 U7315 ( .A1(n4326), .A2(n4325), .ZN(result[3]) );
  NOR2_X4 U7316 ( .A1(net212677), .A2(n4327), .ZN(n4331) );
  NAND2_X2 U7317 ( .A1(n5193), .A2(b[4]), .ZN(n4330) );
  MUX2_X2 U7318 ( .A(n4331), .B(n4330), .S(n4329), .Z(n4375) );
  XNOR2_X2 U7319 ( .A(n4332), .B(net217761), .ZN(n4348) );
  NAND2_X2 U7320 ( .A1(n3998), .A2(a[28]), .ZN(n7067) );
  INV_X4 U7321 ( .A(n7067), .ZN(n4334) );
  INV_X4 U7322 ( .A(a[30]), .ZN(n7889) );
  NOR2_X4 U7323 ( .A1(n4334), .A2(n4333), .ZN(n4336) );
  MUX2_X2 U7324 ( .A(n7817), .B(n7668), .S(net218558), .Z(n4335) );
  NAND2_X2 U7325 ( .A1(n4336), .A2(n4335), .ZN(n7099) );
  NAND2_X2 U7326 ( .A1(n7803), .A2(n7099), .ZN(n4344) );
  NAND2_X2 U7327 ( .A1(net218624), .A2(a[22]), .ZN(n4337) );
  INV_X4 U7328 ( .A(n4337), .ZN(n6645) );
  NOR2_X4 U7329 ( .A1(n3373), .A2(n6645), .ZN(n4339) );
  MUX2_X2 U7330 ( .A(net214224), .B(net213634), .S(net218556), .Z(n4338) );
  NAND2_X2 U7331 ( .A1(n4339), .A2(n4338), .ZN(n4685) );
  NAND2_X2 U7332 ( .A1(n7039), .A2(n4685), .ZN(n4343) );
  NAND2_X2 U7333 ( .A1(net218624), .A2(a[26]), .ZN(n7068) );
  NOR2_X4 U7334 ( .A1(n3332), .A2(n7069), .ZN(n4341) );
  MUX2_X2 U7335 ( .A(net213311), .B(n7816), .S(net218560), .Z(n4340) );
  NAND2_X2 U7336 ( .A1(n4341), .A2(n4340), .ZN(n4947) );
  NAND2_X2 U7337 ( .A1(n7805), .A2(n4947), .ZN(n4342) );
  INV_X4 U7338 ( .A(n6005), .ZN(n4345) );
  NOR2_X4 U7339 ( .A1(n3369), .A2(n4768), .ZN(n4347) );
  AOI211_X2 U7340 ( .C1(n4348), .C2(n3990), .A(n4347), .B(n4346), .ZN(n4374)
         );
  INV_X4 U7341 ( .A(net217654), .ZN(net217736) );
  MUX2_X2 U7342 ( .A(net217736), .B(n4274), .S(net218558), .Z(n4351) );
  NAND2_X2 U7343 ( .A1(n3998), .A2(net219055), .ZN(n4360) );
  NAND2_X2 U7344 ( .A1(net218624), .A2(a[2]), .ZN(n4675) );
  NAND2_X2 U7345 ( .A1(n4360), .A2(n4675), .ZN(n4350) );
  NOR2_X4 U7346 ( .A1(n4351), .A2(n4350), .ZN(n6633) );
  NAND2_X2 U7347 ( .A1(n3998), .A2(a[0]), .ZN(n6632) );
  MUX2_X2 U7348 ( .A(n6633), .B(n6632), .S(net218546), .Z(n7078) );
  NAND2_X2 U7349 ( .A1(n4352), .A2(n3329), .ZN(n4357) );
  INV_X4 U7350 ( .A(n5330), .ZN(n4775) );
  NAND2_X2 U7351 ( .A1(net218624), .A2(a[14]), .ZN(n4353) );
  INV_X4 U7352 ( .A(n4353), .ZN(n5456) );
  NOR2_X4 U7353 ( .A1(n3375), .A2(n5456), .ZN(n4355) );
  MUX2_X2 U7354 ( .A(net216117), .B(net215701), .S(net218560), .Z(n4354) );
  NAND2_X2 U7355 ( .A1(n4355), .A2(n4354), .ZN(n4493) );
  NAND2_X2 U7356 ( .A1(n4775), .A2(n4493), .ZN(n4356) );
  OAI211_X2 U7357 ( .C1(n7078), .C2(n3383), .A(n4357), .B(n4356), .ZN(n4372)
         );
  NAND2_X2 U7358 ( .A1(n4359), .A2(net218556), .ZN(n4763) );
  NAND2_X2 U7359 ( .A1(net218624), .A2(a[6]), .ZN(n4482) );
  NAND4_X2 U7360 ( .A1(n4361), .A2(n4763), .A3(n4482), .A4(n4360), .ZN(n4680)
         );
  INV_X4 U7361 ( .A(n4680), .ZN(n4362) );
  NAND2_X2 U7362 ( .A1(net218624), .A2(a[18]), .ZN(n4363) );
  INV_X4 U7363 ( .A(n4363), .ZN(n6001) );
  NOR2_X4 U7364 ( .A1(n3372), .A2(n6001), .ZN(n4365) );
  MUX2_X2 U7365 ( .A(net215245), .B(net215001), .S(net218558), .Z(n4364) );
  NAND2_X2 U7366 ( .A1(n4365), .A2(n4364), .ZN(n4686) );
  INV_X4 U7367 ( .A(n4686), .ZN(n4950) );
  NAND2_X2 U7368 ( .A1(net218624), .A2(a[10]), .ZN(n4366) );
  INV_X4 U7369 ( .A(n4366), .ZN(n4939) );
  NOR2_X4 U7370 ( .A1(n3374), .A2(n4939), .ZN(n4368) );
  MUX2_X2 U7371 ( .A(net216885), .B(net216517), .S(net218556), .Z(n4367) );
  NAND2_X2 U7372 ( .A1(n4368), .A2(n4367), .ZN(n4369) );
  INV_X4 U7373 ( .A(n4369), .ZN(n4682) );
  OAI22_X2 U7374 ( .A1(n4950), .A2(n3996), .B1(n4682), .B2(n5332), .ZN(n4370)
         );
  NOR3_X4 U7375 ( .A1(n4372), .A2(n4371), .A3(n4370), .ZN(n4373) );
  NAND4_X2 U7376 ( .A1(n4375), .A2(n3394), .A3(n4374), .A4(n4373), .ZN(
        result[4]) );
  NOR2_X4 U7377 ( .A1(b[5]), .A2(a[5]), .ZN(n4392) );
  INV_X4 U7378 ( .A(n4392), .ZN(n4376) );
  NAND2_X2 U7379 ( .A1(n4376), .A2(net217083), .ZN(net217445) );
  NOR2_X4 U7380 ( .A1(n4378), .A2(n4377), .ZN(n4405) );
  NAND2_X2 U7381 ( .A1(n5193), .A2(b[5]), .ZN(n4382) );
  MUX2_X2 U7382 ( .A(n4382), .B(n4381), .S(n4380), .Z(n4404) );
  INV_X4 U7383 ( .A(n4383), .ZN(n5057) );
  OAI22_X2 U7384 ( .A1(n5057), .A2(n3993), .B1(net216692), .B2(n7079), .ZN(
        n4384) );
  INV_X4 U7385 ( .A(n4384), .ZN(n4387) );
  NAND2_X2 U7386 ( .A1(n7803), .A2(n7380), .ZN(n4385) );
  NAND2_X2 U7387 ( .A1(n4387), .A2(n4385), .ZN(n6112) );
  NAND2_X2 U7388 ( .A1(n7803), .A2(n5054), .ZN(n4386) );
  AOI221_X2 U7389 ( .B1(n5051), .B2(n6112), .C1(n4861), .C2(n6113), .A(n4388), 
        .ZN(n4403) );
  INV_X4 U7390 ( .A(n4389), .ZN(n4391) );
  XNOR2_X2 U7391 ( .A(n4391), .B(n4390), .ZN(n4401) );
  NOR2_X4 U7392 ( .A1(n4395), .A2(n4394), .ZN(n4396) );
  NAND2_X2 U7393 ( .A1(n4397), .A2(n4396), .ZN(n4400) );
  NAND2_X2 U7394 ( .A1(n5446), .A2(n7805), .ZN(n7053) );
  NAND2_X2 U7395 ( .A1(n6851), .A2(n6100), .ZN(n4398) );
  AOI211_X2 U7396 ( .C1(n4401), .C2(n3990), .A(n4400), .B(n4399), .ZN(n4402)
         );
  NAND4_X2 U7397 ( .A1(n4405), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(
        result[5]) );
  NOR2_X4 U7398 ( .A1(b[6]), .A2(a[6]), .ZN(n4425) );
  INV_X4 U7399 ( .A(n4425), .ZN(n4406) );
  NAND2_X2 U7400 ( .A1(b[6]), .A2(a[6]), .ZN(net216979) );
  NAND2_X2 U7401 ( .A1(n4406), .A2(net216979), .ZN(n4592) );
  NOR2_X4 U7402 ( .A1(n4408), .A2(n4407), .ZN(n4441) );
  NOR2_X4 U7403 ( .A1(b[6]), .A2(net218659), .ZN(n4409) );
  NAND2_X2 U7404 ( .A1(n5193), .A2(b[6]), .ZN(n4412) );
  MUX2_X2 U7405 ( .A(n4413), .B(n4412), .S(n4411), .Z(n4440) );
  AOI22_X2 U7406 ( .A1(n7039), .A2(n4778), .B1(n7805), .B2(n5178), .ZN(n4417)
         );
  NAND2_X2 U7407 ( .A1(n7803), .A2(n7831), .ZN(n4414) );
  NAND2_X2 U7408 ( .A1(n4417), .A2(n4414), .ZN(n6137) );
  NAND2_X2 U7409 ( .A1(n7803), .A2(n7829), .ZN(n4415) );
  INV_X4 U7410 ( .A(n4418), .ZN(n4419) );
  MUX2_X2 U7411 ( .A(n4484), .B(net217654), .S(net218558), .Z(n4421) );
  NAND2_X2 U7412 ( .A1(n4422), .A2(n4421), .ZN(n5739) );
  INV_X4 U7413 ( .A(n5739), .ZN(n6273) );
  AOI221_X2 U7414 ( .B1(n5051), .B2(n6137), .C1(n4861), .C2(n6131), .A(n4423), 
        .ZN(n4439) );
  XNOR2_X2 U7415 ( .A(n4424), .B(n3354), .ZN(n4437) );
  INV_X4 U7416 ( .A(n4427), .ZN(n4777) );
  INV_X4 U7417 ( .A(n4774), .ZN(n5181) );
  NOR2_X4 U7418 ( .A1(n4429), .A2(n4428), .ZN(n4430) );
  NAND2_X2 U7419 ( .A1(n4431), .A2(n4430), .ZN(n4436) );
  INV_X4 U7420 ( .A(n4432), .ZN(n4434) );
  NAND2_X2 U7421 ( .A1(n6851), .A2(n6272), .ZN(n4433) );
  AOI211_X2 U7422 ( .C1(n4437), .C2(n3990), .A(n4436), .B(n4435), .ZN(n4438)
         );
  NAND4_X2 U7423 ( .A1(n4441), .A2(n4440), .A3(n4439), .A4(n4438), .ZN(
        result[6]) );
  NOR2_X4 U7424 ( .A1(b[7]), .A2(a[7]), .ZN(net217608) );
  INV_X4 U7425 ( .A(net217608), .ZN(net217631) );
  NAND2_X2 U7426 ( .A1(b[7]), .A2(a[7]), .ZN(net216394) );
  NOR2_X4 U7427 ( .A1(n4442), .A2(net217630), .ZN(n4472) );
  NAND2_X2 U7428 ( .A1(n5193), .A2(b[7]), .ZN(n4446) );
  MUX2_X2 U7429 ( .A(n4446), .B(n4445), .S(n4444), .Z(n4471) );
  NAND4_X2 U7430 ( .A1(net217621), .A2(n4449), .A3(n4448), .A4(n4447), .ZN(
        n6451) );
  AOI22_X2 U7431 ( .A1(n3992), .A2(n4865), .B1(n7039), .B2(n4450), .ZN(n4452)
         );
  INV_X4 U7432 ( .A(n6467), .ZN(n4451) );
  NAND2_X2 U7433 ( .A1(n4452), .A2(n6636), .ZN(n6469) );
  INV_X4 U7434 ( .A(n6469), .ZN(n4453) );
  NOR3_X4 U7435 ( .A1(n3205), .A2(n4455), .A3(n4454), .ZN(n4470) );
  INV_X4 U7436 ( .A(n4456), .ZN(n4458) );
  XNOR2_X2 U7437 ( .A(n4458), .B(n4457), .ZN(n4468) );
  NOR2_X4 U7438 ( .A1(n4462), .A2(n4461), .ZN(n4463) );
  NAND2_X2 U7439 ( .A1(n4464), .A2(n4463), .ZN(n4467) );
  NAND2_X2 U7440 ( .A1(n6851), .A2(n5315), .ZN(n4465) );
  AOI211_X2 U7441 ( .C1(n4468), .C2(n3990), .A(n4467), .B(n4466), .ZN(n4469)
         );
  NAND4_X2 U7442 ( .A1(n4472), .A2(n4471), .A3(n4470), .A4(n4469), .ZN(
        result[7]) );
  NOR2_X4 U7443 ( .A1(b[8]), .A2(a[8]), .ZN(n4494) );
  INV_X4 U7444 ( .A(n4494), .ZN(n4473) );
  NAND2_X2 U7445 ( .A1(n4473), .A2(net216097), .ZN(n4607) );
  NOR2_X4 U7446 ( .A1(n4475), .A2(n4474), .ZN(n4502) );
  NOR2_X4 U7447 ( .A1(b[8]), .A2(net218659), .ZN(n4476) );
  NAND2_X2 U7448 ( .A1(n5193), .A2(b[8]), .ZN(n4479) );
  INV_X4 U7449 ( .A(n4477), .ZN(n4478) );
  MUX2_X2 U7450 ( .A(n4480), .B(n4479), .S(n4478), .Z(n4501) );
  XNOR2_X2 U7451 ( .A(n4481), .B(net217584), .ZN(n4491) );
  INV_X4 U7452 ( .A(n4482), .ZN(n4483) );
  NOR2_X4 U7453 ( .A1(n3374), .A2(n4483), .ZN(n4487) );
  MUX2_X2 U7454 ( .A(n4485), .B(n3910), .S(net218556), .Z(n4486) );
  NAND2_X2 U7455 ( .A1(n4487), .A2(n4486), .ZN(n5449) );
  INV_X4 U7456 ( .A(n5449), .ZN(n7081) );
  INV_X4 U7457 ( .A(n7036), .ZN(n6639) );
  NAND2_X2 U7458 ( .A1(n6639), .A2(net218538), .ZN(n4488) );
  AOI211_X2 U7459 ( .C1(n4491), .C2(n3990), .A(n4490), .B(n4489), .ZN(n4500)
         );
  INV_X4 U7460 ( .A(n4685), .ZN(n4949) );
  INV_X4 U7461 ( .A(n6632), .ZN(n5451) );
  NAND2_X2 U7462 ( .A1(n5446), .A2(n7803), .ZN(n6984) );
  INV_X4 U7463 ( .A(n6984), .ZN(n7033) );
  NAND2_X2 U7464 ( .A1(n5451), .A2(n7033), .ZN(n4492) );
  OAI221_X2 U7465 ( .B1(n4949), .B2(n3996), .C1(n4682), .C2(n4942), .A(n4492), 
        .ZN(n4498) );
  INV_X4 U7466 ( .A(n4493), .ZN(n4943) );
  OAI22_X2 U7467 ( .A1(n4943), .A2(n5332), .B1(n4950), .B2(n5330), .ZN(n4497)
         );
  AOI22_X2 U7468 ( .A1(n7039), .A2(n4947), .B1(n7805), .B2(n7099), .ZN(n6652)
         );
  NAND2_X2 U7469 ( .A1(n4860), .A2(n4768), .ZN(n4952) );
  INV_X4 U7470 ( .A(n4952), .ZN(n4495) );
  NOR3_X4 U7471 ( .A1(n4498), .A2(n4497), .A3(n4496), .ZN(n4499) );
  NAND4_X2 U7472 ( .A1(n4502), .A2(n4501), .A3(n4500), .A4(n4499), .ZN(
        result[8]) );
  NAND2_X2 U7473 ( .A1(a[31]), .A2(net212023), .ZN(n4572) );
  NAND2_X2 U7474 ( .A1(net217362), .A2(n4572), .ZN(net217356) );
  INV_X4 U7475 ( .A(net217356), .ZN(net211993) );
  NAND2_X2 U7476 ( .A1(net211993), .A2(a[30]), .ZN(n4574) );
  XNOR2_X2 U7477 ( .A(a[29]), .B(b[29]), .ZN(n7230) );
  XNOR2_X2 U7478 ( .A(a[27]), .B(b[27]), .ZN(n7055) );
  XNOR2_X2 U7479 ( .A(a[25]), .B(b[25]), .ZN(n4647) );
  XNOR2_X2 U7480 ( .A(a[24]), .B(b[24]), .ZN(n4590) );
  INV_X4 U7481 ( .A(n4590), .ZN(n6650) );
  INV_X4 U7482 ( .A(b[23]), .ZN(net214747) );
  NAND2_X2 U7483 ( .A1(a[23]), .A2(net214747), .ZN(n4560) );
  XNOR2_X2 U7484 ( .A(a[20]), .B(b[20]), .ZN(n4504) );
  INV_X4 U7485 ( .A(n4504), .ZN(n5998) );
  NOR2_X4 U7486 ( .A1(n3378), .A2(n5998), .ZN(n4505) );
  XNOR2_X2 U7487 ( .A(a[19]), .B(b[19]), .ZN(n4626) );
  XNOR2_X2 U7488 ( .A(a[21]), .B(b[21]), .ZN(n6108) );
  XNOR2_X2 U7489 ( .A(a[22]), .B(b[22]), .ZN(n6144) );
  NAND4_X2 U7490 ( .A1(n4505), .A2(n4626), .A3(n6108), .A4(n6144), .ZN(n4591)
         );
  INV_X4 U7491 ( .A(n4591), .ZN(n4633) );
  XNOR2_X2 U7492 ( .A(a[16]), .B(b[16]), .ZN(n4623) );
  NOR2_X4 U7493 ( .A1(a[15]), .A2(b[15]), .ZN(n5328) );
  INV_X4 U7494 ( .A(n5328), .ZN(n4506) );
  NAND2_X2 U7495 ( .A1(n4506), .A2(n7589), .ZN(n5190) );
  INV_X4 U7496 ( .A(n5190), .ZN(n4576) );
  NOR2_X4 U7497 ( .A1(b[13]), .A2(a[13]), .ZN(net216698) );
  INV_X4 U7498 ( .A(net216698), .ZN(net217552) );
  INV_X4 U7499 ( .A(net216856), .ZN(net217464) );
  NOR2_X4 U7500 ( .A1(b[11]), .A2(a[11]), .ZN(n4863) );
  INV_X4 U7501 ( .A(n4863), .ZN(n4507) );
  NAND2_X2 U7502 ( .A1(n4507), .A2(n6382), .ZN(n4787) );
  INV_X4 U7503 ( .A(n4787), .ZN(n4534) );
  NOR2_X4 U7504 ( .A1(b[10]), .A2(a[10]), .ZN(net217169) );
  INV_X4 U7505 ( .A(net217169), .ZN(net217550) );
  OAI21_X4 U7506 ( .B1(net215584), .B2(n4508), .A(net217299), .ZN(n4610) );
  INV_X4 U7507 ( .A(n4610), .ZN(n4532) );
  NAND2_X2 U7508 ( .A1(a[2]), .A2(net218554), .ZN(n4513) );
  NAND2_X2 U7509 ( .A1(a[0]), .A2(net218578), .ZN(n4509) );
  INV_X4 U7510 ( .A(net217427), .ZN(net217541) );
  AOI21_X4 U7511 ( .B1(n4513), .B2(n4512), .A(net217541), .ZN(n4519) );
  INV_X4 U7512 ( .A(net217445), .ZN(net217529) );
  INV_X4 U7513 ( .A(net217439), .ZN(net217526) );
  INV_X4 U7514 ( .A(n4607), .ZN(n4514) );
  NOR2_X4 U7515 ( .A1(net217526), .A2(n4514), .ZN(n4515) );
  INV_X4 U7516 ( .A(n4603), .ZN(n4517) );
  OAI21_X4 U7517 ( .B1(n4519), .B2(n4518), .A(n4517), .ZN(n4528) );
  NOR2_X4 U7518 ( .A1(b[5]), .A2(net218456), .ZN(n4521) );
  NOR2_X4 U7519 ( .A1(b[7]), .A2(net218442), .ZN(n4524) );
  NAND2_X2 U7520 ( .A1(a[8]), .A2(net218514), .ZN(n4526) );
  NAND3_X2 U7521 ( .A1(n4528), .A2(n4527), .A3(n4526), .ZN(n4531) );
  NOR2_X4 U7522 ( .A1(b[10]), .A2(net218420), .ZN(n4530) );
  INV_X4 U7523 ( .A(net217299), .ZN(net217517) );
  AOI211_X2 U7524 ( .C1(n4532), .C2(n4531), .A(n4530), .B(n4529), .ZN(n4533)
         );
  OAI21_X4 U7525 ( .B1(n4534), .B2(n4533), .A(net217512), .ZN(n4537) );
  NOR2_X4 U7526 ( .A1(b[12]), .A2(a[12]), .ZN(n4951) );
  INV_X4 U7527 ( .A(n4951), .ZN(n4535) );
  NAND2_X2 U7528 ( .A1(n4535), .A2(net214022), .ZN(n4875) );
  NOR2_X4 U7529 ( .A1(b[12]), .A2(net218406), .ZN(n4536) );
  AOI21_X4 U7530 ( .B1(n4537), .B2(n4875), .A(n4536), .ZN(n4538) );
  OAI21_X4 U7531 ( .B1(net217464), .B2(n4538), .A(net217506), .ZN(n4541) );
  NOR2_X4 U7532 ( .A1(a[14]), .A2(b[14]), .ZN(n5172) );
  INV_X4 U7533 ( .A(n5172), .ZN(n4539) );
  NAND2_X2 U7534 ( .A1(a[14]), .A2(b[14]), .ZN(n7246) );
  NAND2_X2 U7535 ( .A1(n4539), .A2(n7246), .ZN(n5067) );
  NOR2_X4 U7536 ( .A1(b[14]), .A2(net218392), .ZN(n4540) );
  AOI21_X4 U7537 ( .B1(n4541), .B2(n5067), .A(n4540), .ZN(n4543) );
  INV_X4 U7538 ( .A(b[15]), .ZN(net217403) );
  NAND2_X2 U7539 ( .A1(a[15]), .A2(net217403), .ZN(n4542) );
  INV_X4 U7540 ( .A(a[16]), .ZN(net216124) );
  AOI21_X4 U7541 ( .B1(n4623), .B2(n4545), .A(n4544), .ZN(n4547) );
  XNOR2_X2 U7542 ( .A(a[17]), .B(b[17]), .ZN(n4579) );
  INV_X4 U7543 ( .A(n4579), .ZN(n5605) );
  INV_X4 U7544 ( .A(b[17]), .ZN(net217497) );
  NAND2_X2 U7545 ( .A1(a[17]), .A2(net217497), .ZN(n4546) );
  INV_X4 U7546 ( .A(a[22]), .ZN(net214758) );
  INV_X4 U7547 ( .A(b[21]), .ZN(net215232) );
  NAND2_X2 U7548 ( .A1(a[21]), .A2(net215232), .ZN(n4554) );
  INV_X4 U7549 ( .A(a[18]), .ZN(net215709) );
  INV_X4 U7550 ( .A(a[19]), .ZN(net215499) );
  AOI21_X2 U7551 ( .B1(n4549), .B2(n4626), .A(n4548), .ZN(n4550) );
  INV_X4 U7552 ( .A(a[20]), .ZN(net215252) );
  INV_X4 U7553 ( .A(n6144), .ZN(n4635) );
  XNOR2_X2 U7554 ( .A(a[23]), .B(b[23]), .ZN(n6463) );
  NAND2_X2 U7555 ( .A1(n4590), .A2(n6463), .ZN(n4642) );
  INV_X4 U7556 ( .A(b[24]), .ZN(net214247) );
  NAND2_X2 U7557 ( .A1(a[24]), .A2(net214247), .ZN(n4558) );
  OAI221_X2 U7558 ( .B1(n6650), .B2(n4560), .C1(n4559), .C2(n4642), .A(n4558), 
        .ZN(n4562) );
  INV_X4 U7559 ( .A(a[25]), .ZN(net213919) );
  AOI21_X2 U7560 ( .B1(n4647), .B2(n4562), .A(n4561), .ZN(n4565) );
  XNOR2_X2 U7561 ( .A(a[26]), .B(b[26]), .ZN(n4563) );
  INV_X4 U7562 ( .A(n4563), .ZN(n7001) );
  INV_X4 U7563 ( .A(b[26]), .ZN(net217478) );
  NAND2_X2 U7564 ( .A1(a[26]), .A2(net217478), .ZN(n4564) );
  INV_X4 U7565 ( .A(a[27]), .ZN(n7054) );
  AOI21_X4 U7566 ( .B1(n7055), .B2(n4567), .A(n4566), .ZN(n4569) );
  XNOR2_X2 U7567 ( .A(a[28]), .B(b[28]), .ZN(n7089) );
  INV_X4 U7568 ( .A(n7089), .ZN(n4653) );
  INV_X4 U7569 ( .A(b[28]), .ZN(net212989) );
  NAND2_X2 U7570 ( .A1(a[28]), .A2(net212989), .ZN(n4568) );
  INV_X4 U7571 ( .A(a[29]), .ZN(n7387) );
  XNOR2_X2 U7572 ( .A(b[30]), .B(a[30]), .ZN(n7825) );
  NAND2_X2 U7573 ( .A1(net211993), .A2(n7825), .ZN(n4658) );
  OAI221_X2 U7574 ( .B1(b[30]), .B2(n4574), .C1(n4573), .C2(n4658), .A(n4572), 
        .ZN(n4575) );
  XNOR2_X2 U7575 ( .A(n4575), .B(net217356), .ZN(n4664) );
  NAND2_X2 U7576 ( .A1(n4787), .A2(net217427), .ZN(n4577) );
  INV_X4 U7577 ( .A(n4875), .ZN(n4616) );
  INV_X4 U7578 ( .A(n5067), .ZN(n4620) );
  NOR4_X2 U7579 ( .A1(n4577), .A2(n4616), .A3(n4620), .A4(net217464), .ZN(
        n4587) );
  INV_X4 U7580 ( .A(n4647), .ZN(n6859) );
  NAND4_X2 U7581 ( .A1(n4578), .A2(n7055), .A3(n7230), .A4(n7089), .ZN(n4585)
         );
  NAND2_X2 U7582 ( .A1(n4579), .A2(n4623), .ZN(n4584) );
  INV_X4 U7583 ( .A(n4701), .ZN(n4580) );
  NAND2_X2 U7584 ( .A1(n4580), .A2(n4700), .ZN(n4581) );
  NAND3_X2 U7585 ( .A1(net217433), .A2(n4582), .A3(n4581), .ZN(n4583) );
  NAND4_X2 U7586 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4661)
         );
  INV_X4 U7587 ( .A(n4661), .ZN(n4668) );
  NAND2_X2 U7588 ( .A1(n4668), .A2(net217346), .ZN(n4667) );
  NAND2_X2 U7589 ( .A1(n4664), .A2(n4667), .ZN(n4666) );
  NAND2_X2 U7590 ( .A1(b[23]), .A2(n4590), .ZN(n4644) );
  NAND2_X2 U7591 ( .A1(b[9]), .A2(net217299), .ZN(n4612) );
  NAND2_X2 U7592 ( .A1(b[7]), .A2(net218442), .ZN(n4597) );
  NAND2_X2 U7593 ( .A1(b[5]), .A2(net218456), .ZN(n4594) );
  INV_X4 U7594 ( .A(n4592), .ZN(n4593) );
  NAND2_X2 U7595 ( .A1(n4597), .A2(n4596), .ZN(n4608) );
  NOR2_X4 U7596 ( .A1(a[8]), .A2(net218514), .ZN(n4606) );
  NOR2_X4 U7597 ( .A1(a[3]), .A2(net218544), .ZN(n4601) );
  AOI21_X4 U7598 ( .B1(n4602), .B2(net217427), .A(n4601), .ZN(n4604) );
  NOR2_X4 U7599 ( .A1(n4604), .A2(n4603), .ZN(n4605) );
  NAND2_X2 U7600 ( .A1(b[10]), .A2(net218420), .ZN(n4609) );
  OAI221_X2 U7601 ( .B1(a[9]), .B2(n4612), .C1(n4611), .C2(n4610), .A(n4609), 
        .ZN(n4613) );
  AOI21_X2 U7602 ( .B1(n4613), .B2(n4787), .A(net217414), .ZN(n4615) );
  NAND2_X2 U7603 ( .A1(b[12]), .A2(net218406), .ZN(n4614) );
  OAI21_X4 U7604 ( .B1(n4616), .B2(n4615), .A(n4614), .ZN(n4617) );
  AOI21_X4 U7605 ( .B1(n4617), .B2(net216856), .A(net217408), .ZN(n4619) );
  NAND2_X2 U7606 ( .A1(b[14]), .A2(net218392), .ZN(n4618) );
  OAI21_X4 U7607 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n4622) );
  INV_X4 U7608 ( .A(n4623), .ZN(n5453) );
  NAND2_X2 U7609 ( .A1(b[16]), .A2(net216124), .ZN(n4624) );
  INV_X4 U7610 ( .A(n4626), .ZN(n5874) );
  INV_X4 U7611 ( .A(b[18]), .ZN(net217396) );
  NOR2_X4 U7612 ( .A1(n5874), .A2(net217396), .ZN(n4628) );
  INV_X4 U7613 ( .A(b[19]), .ZN(net217395) );
  AOI21_X4 U7614 ( .B1(n4628), .B2(net215709), .A(n4627), .ZN(n4630) );
  NAND2_X2 U7615 ( .A1(b[20]), .A2(net215252), .ZN(n4629) );
  NAND3_X2 U7616 ( .A1(n4633), .A2(b[17]), .A3(net218378), .ZN(n4634) );
  INV_X4 U7617 ( .A(b[22]), .ZN(net214984) );
  INV_X4 U7618 ( .A(a[24]), .ZN(net214219) );
  NAND2_X2 U7619 ( .A1(b[24]), .A2(net214219), .ZN(n4641) );
  OAI221_X2 U7620 ( .B1(a[23]), .B2(n4644), .C1(n4643), .C2(n4642), .A(n4641), 
        .ZN(n4646) );
  INV_X4 U7621 ( .A(b[25]), .ZN(net217376) );
  NOR2_X4 U7622 ( .A1(a[25]), .A2(net217376), .ZN(n4645) );
  AOI21_X2 U7623 ( .B1(n4647), .B2(n4646), .A(n4645), .ZN(n4649) );
  INV_X4 U7624 ( .A(a[26]), .ZN(n6999) );
  NAND2_X2 U7625 ( .A1(b[26]), .A2(n6999), .ZN(n4648) );
  OAI21_X4 U7626 ( .B1(n4649), .B2(n7001), .A(n4648), .ZN(n4651) );
  INV_X4 U7627 ( .A(b[27]), .ZN(net213272) );
  NOR2_X4 U7628 ( .A1(a[27]), .A2(net213272), .ZN(n4650) );
  AOI21_X4 U7629 ( .B1(n7055), .B2(n4651), .A(n4650), .ZN(n4654) );
  INV_X4 U7630 ( .A(a[28]), .ZN(n7206) );
  NAND2_X2 U7631 ( .A1(b[28]), .A2(n7206), .ZN(n4652) );
  OAI21_X4 U7632 ( .B1(n4654), .B2(n4653), .A(n4652), .ZN(n4656) );
  INV_X4 U7633 ( .A(b[29]), .ZN(net217365) );
  NOR2_X4 U7634 ( .A1(a[29]), .A2(net217365), .ZN(n4655) );
  AOI21_X4 U7635 ( .B1(n7230), .B2(n4656), .A(n4655), .ZN(n4659) );
  INV_X4 U7636 ( .A(net217362), .ZN(net217361) );
  AOI21_X4 U7637 ( .B1(net217360), .B2(n7889), .A(net217361), .ZN(n4657) );
  OAI21_X4 U7638 ( .B1(n4659), .B2(n4658), .A(n4657), .ZN(n4660) );
  XNOR2_X2 U7639 ( .A(n4660), .B(net217356), .ZN(n4662) );
  NAND2_X2 U7640 ( .A1(n4662), .A2(n4661), .ZN(n4663) );
  MUX2_X2 U7641 ( .A(n4664), .B(n4663), .S(op[0]), .Z(n4665) );
  MUX2_X2 U7642 ( .A(n4666), .B(n4665), .S(op[1]), .Z(net217348) );
  INV_X4 U7643 ( .A(n4667), .ZN(n4670) );
  OAI21_X4 U7644 ( .B1(n4670), .B2(n4669), .A(net217344), .ZN(n4671) );
  MUX2_X2 U7645 ( .A(net217340), .B(n4671), .S(op[2]), .Z(n4708) );
  NAND2_X2 U7646 ( .A1(n4673), .A2(n4672), .ZN(n4706) );
  NAND2_X2 U7647 ( .A1(n4674), .A2(a[3]), .ZN(n4676) );
  NAND2_X2 U7648 ( .A1(n4676), .A2(n4675), .ZN(n4679) );
  NAND2_X2 U7649 ( .A1(n6632), .A2(n4677), .ZN(n4678) );
  NAND2_X2 U7650 ( .A1(n7039), .A2(net218530), .ZN(n7818) );
  INV_X4 U7651 ( .A(n7818), .ZN(n7866) );
  NAND2_X2 U7652 ( .A1(n7805), .A2(n4680), .ZN(n4681) );
  NOR2_X4 U7653 ( .A1(n4684), .A2(n4683), .ZN(n4692) );
  NAND2_X2 U7654 ( .A1(n7803), .A2(n4947), .ZN(n4690) );
  NAND2_X2 U7655 ( .A1(n7805), .A2(n4685), .ZN(n4689) );
  NAND2_X2 U7656 ( .A1(n7039), .A2(n4686), .ZN(n4688) );
  NAND2_X2 U7657 ( .A1(n7807), .A2(n7099), .ZN(n4687) );
  NAND4_X2 U7658 ( .A1(n4690), .A2(n4689), .A3(n4688), .A4(n4687), .ZN(n4691)
         );
  INV_X4 U7659 ( .A(n4691), .ZN(n5455) );
  MUX2_X2 U7660 ( .A(n4692), .B(n5455), .S(b[4]), .Z(n4693) );
  NAND2_X2 U7661 ( .A1(n4694), .A2(n4693), .ZN(n4705) );
  NAND2_X2 U7662 ( .A1(n5451), .A2(n7050), .ZN(n4699) );
  NAND2_X2 U7663 ( .A1(n4695), .A2(n4001), .ZN(n4696) );
  NAND3_X2 U7664 ( .A1(n4697), .A2(n3990), .A3(n4696), .ZN(n4698) );
  NAND2_X2 U7665 ( .A1(n4699), .A2(n4698), .ZN(n4704) );
  NAND2_X2 U7666 ( .A1(net218639), .A2(n4700), .ZN(n4702) );
  AOI211_X4 U7667 ( .C1(n4706), .C2(n4705), .A(n4704), .B(n4703), .ZN(n4707)
         );
  NAND3_X2 U7668 ( .A1(n4709), .A2(n4708), .A3(n4707), .ZN(result[0]) );
  NOR2_X4 U7669 ( .A1(n4710), .A2(net217298), .ZN(n4786) );
  NAND2_X2 U7670 ( .A1(n5193), .A2(b[10]), .ZN(n4758) );
  NAND2_X2 U7671 ( .A1(b[6]), .A2(net219055), .ZN(n4727) );
  INV_X4 U7672 ( .A(n4727), .ZN(n4726) );
  NAND2_X2 U7673 ( .A1(net217282), .A2(net217283), .ZN(n4889) );
  NAND2_X2 U7674 ( .A1(net217273), .A2(net217274), .ZN(n4713) );
  INV_X4 U7675 ( .A(n5044), .ZN(n4712) );
  XNOR2_X2 U7676 ( .A(n4713), .B(net241372), .ZN(net217264) );
  INV_X4 U7677 ( .A(net217264), .ZN(net217267) );
  NAND3_X2 U7678 ( .A1(a[8]), .A2(net217264), .A3(net218548), .ZN(n4799) );
  NAND2_X2 U7679 ( .A1(net216811), .A2(n4799), .ZN(n4717) );
  XOR2_X2 U7680 ( .A(n4717), .B(n4986), .Z(n4715) );
  NAND2_X2 U7681 ( .A1(net218538), .A2(a[7]), .ZN(n4716) );
  INV_X4 U7682 ( .A(n4716), .ZN(n4719) );
  XNOR2_X2 U7683 ( .A(n4721), .B(n4720), .ZN(n4812) );
  INV_X4 U7684 ( .A(n4812), .ZN(n4722) );
  NAND2_X2 U7685 ( .A1(b[4]), .A2(a[6]), .ZN(n4723) );
  INV_X4 U7686 ( .A(n4723), .ZN(n4813) );
  NAND2_X2 U7687 ( .A1(n4813), .A2(n4812), .ZN(net216945) );
  NAND2_X2 U7688 ( .A1(n4815), .A2(n4906), .ZN(n4724) );
  INV_X4 U7689 ( .A(net217240), .ZN(net217238) );
  INV_X4 U7690 ( .A(n4728), .ZN(n4725) );
  AOI21_X4 U7691 ( .B1(n4731), .B2(n4795), .A(n4796), .ZN(n4732) );
  XNOR2_X2 U7692 ( .A(n4733), .B(n4732), .ZN(n4734) );
  INV_X4 U7693 ( .A(n4735), .ZN(n4743) );
  OAI21_X4 U7694 ( .B1(n4743), .B2(n4742), .A(n4741), .ZN(n4881) );
  XNOR2_X2 U7695 ( .A(n4791), .B(n4881), .ZN(n4746) );
  INV_X4 U7696 ( .A(n4746), .ZN(n4744) );
  NAND2_X2 U7697 ( .A1(b[8]), .A2(a[2]), .ZN(n4745) );
  INV_X4 U7698 ( .A(n4745), .ZN(n4747) );
  NAND2_X2 U7699 ( .A1(n4747), .A2(n4746), .ZN(n4829) );
  INV_X4 U7700 ( .A(n4827), .ZN(n4748) );
  XNOR2_X2 U7701 ( .A(n4750), .B(n4749), .ZN(n4752) );
  NAND2_X2 U7702 ( .A1(b[9]), .A2(a[1]), .ZN(n4751) );
  INV_X4 U7703 ( .A(n4751), .ZN(n4753) );
  NAND3_X4 U7704 ( .A1(b[9]), .A2(a[0]), .A3(n4754), .ZN(n4836) );
  XNOR2_X2 U7705 ( .A(n4755), .B(n4836), .ZN(n4756) );
  INV_X4 U7706 ( .A(n4756), .ZN(n4845) );
  MUX2_X2 U7707 ( .A(n4758), .B(n4757), .S(n4845), .Z(n4785) );
  XNOR2_X2 U7708 ( .A(n4000), .B(b[10]), .ZN(n4850) );
  XNOR2_X2 U7709 ( .A(n4850), .B(net218420), .ZN(n4849) );
  OAI22_X2 U7710 ( .A1(n4761), .A2(net218428), .B1(n4760), .B2(n4759), .ZN(
        n4853) );
  XNOR2_X2 U7711 ( .A(n4849), .B(n4853), .ZN(n4771) );
  INV_X4 U7712 ( .A(n7829), .ZN(n4762) );
  NAND2_X2 U7713 ( .A1(n7039), .A2(n5178), .ZN(n4772) );
  OAI211_X2 U7714 ( .C1(n4762), .C2(n3993), .A(n4772), .B(n6636), .ZN(n6995)
         );
  INV_X4 U7715 ( .A(n6995), .ZN(n4769) );
  INV_X4 U7716 ( .A(n6272), .ZN(n4766) );
  NAND4_X2 U7717 ( .A1(net217179), .A2(n4764), .A3(n4763), .A4(net217182), 
        .ZN(n6278) );
  NAND2_X2 U7718 ( .A1(n7039), .A2(n6278), .ZN(n4765) );
  OAI221_X2 U7719 ( .B1(n4766), .B2(n3995), .C1(n6273), .C2(n3993), .A(n4765), 
        .ZN(n7000) );
  NAND2_X2 U7720 ( .A1(n5446), .A2(n7000), .ZN(n4767) );
  AOI21_X2 U7721 ( .B1(n4771), .B2(n3990), .A(n4770), .ZN(n4784) );
  INV_X4 U7722 ( .A(n4772), .ZN(n4773) );
  NAND2_X2 U7723 ( .A1(n4775), .A2(n4774), .ZN(n4776) );
  OAI211_X2 U7724 ( .C1(n6977), .C2(n4860), .A(n3410), .B(n4776), .ZN(n4782)
         );
  INV_X4 U7725 ( .A(n4778), .ZN(n5180) );
  OAI22_X2 U7726 ( .A1(n5180), .A2(n3996), .B1(n4779), .B2(n5332), .ZN(n4780)
         );
  NOR3_X2 U7727 ( .A1(n4782), .A2(n4781), .A3(n4780), .ZN(n4783) );
  NAND4_X2 U7728 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), .ZN(
        result[10]) );
  NOR2_X4 U7729 ( .A1(n4789), .A2(n4788), .ZN(n4874) );
  NAND2_X2 U7730 ( .A1(n5193), .A2(b[11]), .ZN(n4848) );
  OAI211_X2 U7731 ( .C1(n4796), .C2(n4731), .A(n4795), .B(n4794), .ZN(n4886)
         );
  NAND2_X2 U7732 ( .A1(b[5]), .A2(a[6]), .ZN(net217088) );
  NAND2_X2 U7733 ( .A1(b[4]), .A2(a[7]), .ZN(n4810) );
  INV_X4 U7734 ( .A(n4810), .ZN(n4809) );
  NAND2_X2 U7735 ( .A1(net218558), .A2(a[10]), .ZN(net216968) );
  INV_X4 U7736 ( .A(net217121), .ZN(net217122) );
  NAND3_X4 U7737 ( .A1(net217122), .A2(a[9]), .A3(net218546), .ZN(n4893) );
  INV_X4 U7738 ( .A(n4893), .ZN(n4987) );
  NAND2_X2 U7739 ( .A1(net218548), .A2(a[9]), .ZN(n4797) );
  NAND2_X2 U7740 ( .A1(n4797), .A2(net217121), .ZN(n4988) );
  NAND2_X2 U7741 ( .A1(net217118), .A2(n4798), .ZN(n4800) );
  INV_X4 U7742 ( .A(n4799), .ZN(n4989) );
  NAND2_X2 U7743 ( .A1(net218538), .A2(a[8]), .ZN(n4802) );
  NAND2_X2 U7744 ( .A1(n3775), .A2(n4802), .ZN(n4892) );
  INV_X4 U7745 ( .A(n4802), .ZN(n4804) );
  NAND2_X2 U7746 ( .A1(n4892), .A2(n4981), .ZN(n4807) );
  NAND3_X4 U7747 ( .A1(n3782), .A2(net219368), .A3(net218072), .ZN(n4887) );
  NAND2_X2 U7748 ( .A1(b[6]), .A2(a[5]), .ZN(n4817) );
  INV_X4 U7749 ( .A(n4817), .ZN(n4818) );
  XNOR2_X2 U7750 ( .A(n4883), .B(n4819), .ZN(net217070) );
  INV_X4 U7751 ( .A(net217070), .ZN(net217072) );
  NAND2_X2 U7752 ( .A1(b[7]), .A2(net219055), .ZN(net217071) );
  XNOR2_X2 U7753 ( .A(n4820), .B(net217069), .ZN(n4822) );
  INV_X4 U7754 ( .A(n4822), .ZN(n4821) );
  OAI21_X4 U7755 ( .B1(net218470), .B2(net218514), .A(n4821), .ZN(n5009) );
  NAND3_X2 U7756 ( .A1(a[3]), .A2(n4822), .A3(b[8]), .ZN(n5080) );
  NAND2_X2 U7757 ( .A1(n5009), .A2(n5080), .ZN(n4920) );
  INV_X4 U7758 ( .A(n4920), .ZN(n4833) );
  INV_X4 U7759 ( .A(n4823), .ZN(n4831) );
  INV_X4 U7760 ( .A(n4824), .ZN(n4828) );
  INV_X4 U7761 ( .A(n4825), .ZN(n4826) );
  AOI21_X4 U7762 ( .B1(n4828), .B2(n4827), .A(n4826), .ZN(n4830) );
  OAI21_X4 U7763 ( .B1(n4831), .B2(n4830), .A(n4829), .ZN(n5008) );
  XNOR2_X2 U7764 ( .A(n4832), .B(n4833), .ZN(n5020) );
  INV_X4 U7765 ( .A(n4834), .ZN(n4837) );
  OAI21_X4 U7766 ( .B1(n4837), .B2(n4836), .A(n4835), .ZN(n5019) );
  INV_X4 U7767 ( .A(n5019), .ZN(n4839) );
  NAND2_X2 U7768 ( .A1(b[10]), .A2(a[1]), .ZN(n4843) );
  INV_X4 U7769 ( .A(n4843), .ZN(n4929) );
  INV_X4 U7770 ( .A(n4844), .ZN(n4841) );
  INV_X4 U7771 ( .A(n4965), .ZN(n4842) );
  NAND3_X4 U7772 ( .A1(b[10]), .A2(a[0]), .A3(n4845), .ZN(n4928) );
  XNOR2_X2 U7773 ( .A(n4846), .B(n4928), .ZN(n4934) );
  MUX2_X2 U7774 ( .A(n4848), .B(n4847), .S(n4934), .Z(n4873) );
  INV_X4 U7775 ( .A(n4849), .ZN(n4852) );
  INV_X4 U7776 ( .A(n4850), .ZN(n4851) );
  AOI22_X2 U7777 ( .A1(n4853), .A2(n4852), .B1(a[10]), .B2(n4851), .ZN(
        net217000) );
  XNOR2_X2 U7778 ( .A(n4000), .B(b[11]), .ZN(net216998) );
  INV_X4 U7779 ( .A(net217001), .ZN(net217031) );
  XNOR2_X2 U7780 ( .A(net217000), .B(net217031), .ZN(n4859) );
  NAND2_X2 U7781 ( .A1(n7805), .A2(n6451), .ZN(n4854) );
  OAI221_X2 U7782 ( .B1(net214476), .B2(n7079), .C1(n6453), .C2(n3995), .A(
        n4854), .ZN(n4855) );
  INV_X4 U7783 ( .A(n4855), .ZN(n7059) );
  INV_X4 U7784 ( .A(n4942), .ZN(n5321) );
  NAND2_X2 U7785 ( .A1(n5321), .A2(n4856), .ZN(n4857) );
  AOI21_X2 U7786 ( .B1(n4859), .B2(n3990), .A(n4858), .ZN(n4872) );
  NAND2_X2 U7787 ( .A1(n6639), .A2(n7079), .ZN(n5176) );
  NAND2_X2 U7788 ( .A1(n4861), .A2(n7039), .ZN(n4862) );
  INV_X4 U7789 ( .A(n4862), .ZN(n5174) );
  OAI211_X2 U7790 ( .C1(n7038), .C2(n3393), .A(n5176), .B(n4866), .ZN(n4870)
         );
  OAI22_X2 U7791 ( .A1(n4867), .A2(n5332), .B1(net216306), .B2(n5330), .ZN(
        n4868) );
  NOR3_X4 U7792 ( .A1(n4870), .A2(n4869), .A3(n4868), .ZN(n4871) );
  NAND4_X2 U7793 ( .A1(n4874), .A2(n4873), .A3(n4872), .A4(n4871), .ZN(
        result[11]) );
  XNOR2_X2 U7794 ( .A(n4000), .B(b[12]), .ZN(n5039) );
  XNOR2_X2 U7795 ( .A(n5039), .B(net218406), .ZN(n5038) );
  XNOR2_X2 U7796 ( .A(n5038), .B(net216716), .ZN(n4877) );
  AOI21_X2 U7797 ( .B1(n4877), .B2(n3990), .A(n4876), .ZN(n4960) );
  NAND2_X2 U7798 ( .A1(n5193), .A2(b[12]), .ZN(n4938) );
  INV_X4 U7799 ( .A(n5009), .ZN(n4879) );
  XNOR2_X2 U7800 ( .A(n4819), .B(n4883), .ZN(net216987) );
  NAND2_X2 U7801 ( .A1(n4884), .A2(net216839), .ZN(n4910) );
  AOI21_X2 U7802 ( .B1(n4986), .B2(net216811), .A(n4989), .ZN(n4894) );
  NAND2_X2 U7803 ( .A1(net218548), .A2(a[10]), .ZN(n4896) );
  INV_X4 U7804 ( .A(net216958), .ZN(net216960) );
  XNOR2_X2 U7805 ( .A(n4898), .B(n5098), .ZN(n4901) );
  NAND2_X2 U7806 ( .A1(net218538), .A2(a[9]), .ZN(n4900) );
  INV_X4 U7807 ( .A(n4900), .ZN(n4902) );
  XNOR2_X2 U7808 ( .A(n4904), .B(n4903), .ZN(n4905) );
  INV_X4 U7809 ( .A(net216947), .ZN(net216943) );
  OAI211_X2 U7810 ( .C1(net216943), .C2(net216944), .A(n4906), .B(net223932), 
        .ZN(n4977) );
  XNOR2_X2 U7811 ( .A(n4908), .B(n4909), .ZN(net216936) );
  INV_X4 U7812 ( .A(net219328), .ZN(net216935) );
  NAND2_X2 U7813 ( .A1(b[7]), .A2(a[5]), .ZN(net216929) );
  XNOR2_X2 U7814 ( .A(n4910), .B(net216925), .ZN(n4912) );
  NAND2_X2 U7815 ( .A1(b[8]), .A2(net219055), .ZN(n4911) );
  NAND2_X2 U7816 ( .A1(n4911), .A2(n4912), .ZN(n5083) );
  INV_X4 U7817 ( .A(n4911), .ZN(n4914) );
  INV_X4 U7818 ( .A(n4912), .ZN(n4913) );
  NAND2_X2 U7819 ( .A1(n5083), .A2(n5079), .ZN(n4915) );
  XNOR2_X2 U7820 ( .A(n4916), .B(n4915), .ZN(n4918) );
  NAND2_X2 U7821 ( .A1(a[3]), .A2(b[9]), .ZN(n4917) );
  INV_X4 U7822 ( .A(n4917), .ZN(n4919) );
  NAND2_X2 U7823 ( .A1(n3350), .A2(n4921), .ZN(n5074) );
  XNOR2_X2 U7824 ( .A(n4923), .B(n4922), .ZN(n4926) );
  INV_X4 U7825 ( .A(n4926), .ZN(n4924) );
  NAND2_X2 U7826 ( .A1(b[10]), .A2(a[2]), .ZN(n4925) );
  INV_X4 U7827 ( .A(n4925), .ZN(n4927) );
  NAND2_X2 U7828 ( .A1(n4963), .A2(n4968), .ZN(n4932) );
  INV_X4 U7829 ( .A(n4928), .ZN(n4931) );
  NAND2_X2 U7830 ( .A1(n4931), .A2(n4929), .ZN(n4966) );
  NAND2_X2 U7831 ( .A1(n4931), .A2(n4930), .ZN(n4964) );
  NAND2_X2 U7832 ( .A1(n5290), .A2(n5289), .ZN(n4935) );
  XNOR2_X2 U7833 ( .A(n4935), .B(n5288), .ZN(n4936) );
  INV_X4 U7834 ( .A(n4936), .ZN(n5033) );
  MUX2_X2 U7835 ( .A(n4938), .B(n4937), .S(n5033), .Z(n4959) );
  NOR2_X4 U7836 ( .A1(n3375), .A2(n4939), .ZN(n4941) );
  MUX2_X2 U7837 ( .A(net216517), .B(net216885), .S(net218558), .Z(n4940) );
  NAND2_X2 U7838 ( .A1(n4941), .A2(n4940), .ZN(n5459) );
  INV_X4 U7839 ( .A(n5459), .ZN(n7080) );
  NOR3_X4 U7840 ( .A1(n4946), .A2(n4945), .A3(n4944), .ZN(n4958) );
  INV_X4 U7841 ( .A(n4947), .ZN(n4948) );
  OAI222_X2 U7842 ( .A1(n4950), .A2(n5332), .B1(n4949), .B2(n5330), .C1(n4948), 
        .C2(n3996), .ZN(n4956) );
  NAND3_X2 U7843 ( .A1(n7039), .A2(n7099), .A3(n4952), .ZN(n4953) );
  NAND2_X2 U7844 ( .A1(n4953), .A2(n5176), .ZN(n4954) );
  NOR3_X4 U7845 ( .A1(n4956), .A2(n4955), .A3(n4954), .ZN(n4957) );
  NAND4_X2 U7846 ( .A1(n4960), .A2(n4959), .A3(n4958), .A4(n4957), .ZN(
        result[12]) );
  NOR2_X4 U7847 ( .A1(n4961), .A2(net216855), .ZN(n5066) );
  NAND2_X2 U7848 ( .A1(n5193), .A2(b[13]), .ZN(n5037) );
  NAND2_X2 U7849 ( .A1(b[11]), .A2(a[2]), .ZN(n5137) );
  NAND3_X2 U7850 ( .A1(n4966), .A2(n4965), .A3(n4964), .ZN(n4967) );
  INV_X4 U7851 ( .A(n4967), .ZN(n4969) );
  XNOR2_X2 U7852 ( .A(n5137), .B(n3770), .ZN(n5026) );
  NAND2_X2 U7853 ( .A1(b[9]), .A2(net219055), .ZN(n5016) );
  INV_X4 U7854 ( .A(n5016), .ZN(n5014) );
  NAND2_X2 U7855 ( .A1(b[8]), .A2(a[5]), .ZN(n5005) );
  INV_X4 U7856 ( .A(n5005), .ZN(n5004) );
  NAND2_X2 U7857 ( .A1(net216842), .A2(net216843), .ZN(net216579) );
  NAND2_X2 U7858 ( .A1(b[7]), .A2(a[6]), .ZN(net216761) );
  INV_X4 U7859 ( .A(n4971), .ZN(n4974) );
  NOR2_X4 U7860 ( .A1(n4974), .A2(n4973), .ZN(n4976) );
  OAI21_X4 U7861 ( .B1(n4976), .B2(n3339), .A(n4975), .ZN(n5087) );
  NAND4_X2 U7862 ( .A1(n4979), .A2(n4977), .A3(net216819), .A4(n4978), .ZN(
        n5085) );
  NAND2_X2 U7863 ( .A1(n4980), .A2(n5085), .ZN(net216782) );
  NAND2_X2 U7864 ( .A1(b[4]), .A2(a[9]), .ZN(n4999) );
  OAI21_X4 U7865 ( .B1(n4984), .B2(n4985), .A(n4983), .ZN(n5093) );
  NAND2_X2 U7866 ( .A1(net216811), .A2(n4988), .ZN(n4991) );
  AOI21_X4 U7867 ( .B1(n4989), .B2(n4988), .A(n4987), .ZN(n4990) );
  OAI21_X4 U7868 ( .B1(n4992), .B2(n4991), .A(n4990), .ZN(n4993) );
  INV_X4 U7869 ( .A(n4993), .ZN(n5103) );
  NAND2_X2 U7870 ( .A1(net218558), .A2(a[12]), .ZN(net216632) );
  NAND3_X4 U7871 ( .A1(net216795), .A2(a[11]), .A3(net218546), .ZN(n5101) );
  NAND2_X2 U7872 ( .A1(net218548), .A2(a[11]), .ZN(n4994) );
  NAND2_X2 U7873 ( .A1(n5101), .A2(n5099), .ZN(n4995) );
  XNOR2_X2 U7874 ( .A(n4996), .B(n4995), .ZN(n5089) );
  INV_X4 U7875 ( .A(n3968), .ZN(n4998) );
  NAND2_X2 U7876 ( .A1(net218538), .A2(a[10]), .ZN(n4997) );
  INV_X4 U7877 ( .A(n4997), .ZN(n5090) );
  INV_X4 U7878 ( .A(n4999), .ZN(n5001) );
  XNOR2_X2 U7879 ( .A(net216782), .B(net216783), .ZN(n5002) );
  NAND2_X2 U7880 ( .A1(n5006), .A2(n5005), .ZN(n5082) );
  NOR2_X4 U7881 ( .A1(n5218), .A2(n5007), .ZN(n5013) );
  NAND2_X2 U7882 ( .A1(n5009), .A2(n5008), .ZN(n5078) );
  AOI21_X2 U7883 ( .B1(n5011), .B2(n5083), .A(n5010), .ZN(n5012) );
  XNOR2_X2 U7884 ( .A(n5013), .B(n5012), .ZN(n5015) );
  INV_X4 U7885 ( .A(n5015), .ZN(n5017) );
  INV_X4 U7886 ( .A(n5073), .ZN(n5021) );
  NAND2_X2 U7887 ( .A1(a[3]), .A2(b[10]), .ZN(n5023) );
  NAND2_X2 U7888 ( .A1(n3903), .A2(n5023), .ZN(n5208) );
  INV_X4 U7889 ( .A(n5023), .ZN(n5025) );
  XNOR2_X2 U7890 ( .A(n5026), .B(n5138), .ZN(n5287) );
  INV_X4 U7891 ( .A(n5290), .ZN(n5027) );
  OAI21_X4 U7892 ( .B1(n5027), .B2(n3422), .A(n5289), .ZN(n5028) );
  NAND2_X2 U7893 ( .A1(n5028), .A2(n5287), .ZN(n5141) );
  NAND2_X2 U7894 ( .A1(b[12]), .A2(a[1]), .ZN(n5029) );
  NAND2_X2 U7895 ( .A1(n5030), .A2(n5029), .ZN(n5148) );
  INV_X4 U7896 ( .A(n5029), .ZN(n5032) );
  NAND2_X2 U7897 ( .A1(n5032), .A2(n5031), .ZN(n5149) );
  XNOR2_X2 U7898 ( .A(n5034), .B(n5150), .ZN(n5035) );
  INV_X4 U7899 ( .A(n5035), .ZN(n5157) );
  MUX2_X2 U7900 ( .A(n5037), .B(n5036), .S(n5157), .Z(n5065) );
  INV_X4 U7901 ( .A(n5038), .ZN(n5041) );
  INV_X4 U7902 ( .A(n5039), .ZN(n5040) );
  AOI22_X2 U7903 ( .A1(net216716), .A2(n5041), .B1(a[12]), .B2(n5040), .ZN(
        net216522) );
  XNOR2_X2 U7904 ( .A(n4000), .B(b[13]), .ZN(net216520) );
  INV_X4 U7905 ( .A(net216523), .ZN(net216714) );
  XNOR2_X2 U7906 ( .A(net216522), .B(net216714), .ZN(n5050) );
  INV_X4 U7907 ( .A(n6100), .ZN(n5042) );
  AOI22_X2 U7908 ( .A1(n7039), .A2(n6850), .B1(n7805), .B2(n6123), .ZN(n5046)
         );
  NAND2_X2 U7909 ( .A1(n5321), .A2(net216704), .ZN(n5048) );
  AOI21_X2 U7910 ( .B1(n5050), .B2(n3990), .A(n5049), .ZN(n5064) );
  NAND2_X2 U7911 ( .A1(n5051), .A2(n7039), .ZN(n5052) );
  INV_X4 U7912 ( .A(n5052), .ZN(n5327) );
  NAND2_X2 U7913 ( .A1(n5327), .A2(n7380), .ZN(n5056) );
  NAND3_X2 U7914 ( .A1(n5056), .A2(n5176), .A3(n5055), .ZN(n5062) );
  NOR4_X2 U7915 ( .A1(n5062), .A2(n5061), .A3(n5060), .A4(n5059), .ZN(n5063)
         );
  NAND4_X2 U7916 ( .A1(n5066), .A2(n5065), .A3(n5064), .A4(n5063), .ZN(
        result[13]) );
  NOR2_X4 U7917 ( .A1(n5069), .A2(n5068), .ZN(n5189) );
  NAND2_X2 U7918 ( .A1(n5193), .A2(b[14]), .ZN(n5161) );
  INV_X4 U7919 ( .A(n5208), .ZN(n5072) );
  OAI21_X4 U7920 ( .B1(n5072), .B2(n5071), .A(n5212), .ZN(n5132) );
  NAND3_X2 U7921 ( .A1(n5074), .A2(n5073), .A3(n4840), .ZN(n5075) );
  NAND3_X2 U7922 ( .A1(n3791), .A2(n5076), .A3(n5075), .ZN(n5214) );
  NAND3_X2 U7923 ( .A1(n5081), .A2(n5082), .A3(n5083), .ZN(n5215) );
  INV_X4 U7924 ( .A(n5085), .ZN(n5088) );
  OAI21_X4 U7925 ( .B1(n5088), .B2(n5087), .A(n5086), .ZN(n5223) );
  NAND2_X2 U7926 ( .A1(n5091), .A2(n5360), .ZN(n5095) );
  NAND3_X2 U7927 ( .A1(n5093), .A2(n5092), .A3(n5360), .ZN(n5094) );
  NAND2_X2 U7928 ( .A1(n5095), .A2(n5094), .ZN(n5110) );
  NAND2_X2 U7929 ( .A1(net218536), .A2(a[11]), .ZN(n5107) );
  NAND2_X2 U7930 ( .A1(net218548), .A2(a[12]), .ZN(n5096) );
  INV_X4 U7931 ( .A(net216620), .ZN(net216622) );
  NAND2_X2 U7932 ( .A1(n5096), .A2(net216622), .ZN(n5097) );
  NAND3_X2 U7933 ( .A1(a[12]), .A2(net216620), .A3(net218548), .ZN(n5232) );
  INV_X4 U7934 ( .A(n5099), .ZN(n5105) );
  INV_X4 U7935 ( .A(n5098), .ZN(n5100) );
  XNOR2_X2 U7936 ( .A(n5231), .B(n5233), .ZN(n5108) );
  INV_X4 U7937 ( .A(n5108), .ZN(n5106) );
  INV_X4 U7938 ( .A(n5107), .ZN(n5109) );
  NAND2_X2 U7939 ( .A1(n5109), .A2(n5108), .ZN(n5359) );
  NAND2_X2 U7940 ( .A1(n5246), .A2(n5359), .ZN(n5363) );
  XNOR2_X2 U7941 ( .A(n5110), .B(n5363), .ZN(n5112) );
  NAND2_X2 U7942 ( .A1(b[4]), .A2(a[10]), .ZN(n5111) );
  INV_X4 U7943 ( .A(n5111), .ZN(n5114) );
  INV_X4 U7944 ( .A(n5112), .ZN(n5113) );
  XNOR2_X2 U7945 ( .A(n5116), .B(n5224), .ZN(n5117) );
  OAI21_X4 U7946 ( .B1(n3912), .B2(n3312), .A(net216284), .ZN(n5351) );
  XNOR2_X2 U7947 ( .A(n5118), .B(n5351), .ZN(n5121) );
  NAND2_X2 U7948 ( .A1(b[6]), .A2(a[8]), .ZN(n5120) );
  INV_X4 U7949 ( .A(n5120), .ZN(n5122) );
  INV_X4 U7950 ( .A(net216565), .ZN(net216569) );
  NAND2_X2 U7951 ( .A1(b[8]), .A2(a[6]), .ZN(net216567) );
  OAI21_X4 U7952 ( .B1(net216568), .B2(net216569), .A(net216567), .ZN(n5216)
         );
  INV_X4 U7953 ( .A(net216567), .ZN(net216566) );
  XNOR2_X2 U7954 ( .A(n5125), .B(n5124), .ZN(n5127) );
  NAND2_X2 U7955 ( .A1(b[9]), .A2(a[5]), .ZN(n5126) );
  INV_X4 U7956 ( .A(n5126), .ZN(n5128) );
  XNOR2_X2 U7957 ( .A(n5349), .B(n5129), .ZN(n5205) );
  INV_X4 U7958 ( .A(n5205), .ZN(n5130) );
  XNOR2_X2 U7959 ( .A(n5131), .B(n5132), .ZN(n5135) );
  NAND2_X2 U7960 ( .A1(a[3]), .A2(b[11]), .ZN(n5134) );
  INV_X4 U7961 ( .A(n5134), .ZN(n5136) );
  INV_X4 U7962 ( .A(n5137), .ZN(n5140) );
  XNOR2_X2 U7963 ( .A(n5143), .B(n5142), .ZN(n5146) );
  NAND2_X2 U7964 ( .A1(b[12]), .A2(a[2]), .ZN(n5145) );
  INV_X4 U7965 ( .A(n5145), .ZN(n5147) );
  NAND2_X2 U7966 ( .A1(n5147), .A2(n3419), .ZN(n5201) );
  NAND2_X2 U7967 ( .A1(n5200), .A2(n5201), .ZN(n5152) );
  INV_X4 U7968 ( .A(n5148), .ZN(n5151) );
  OAI21_X4 U7969 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n5199) );
  XNOR2_X2 U7970 ( .A(n5152), .B(n5199), .ZN(n5155) );
  INV_X4 U7971 ( .A(n5155), .ZN(n5153) );
  NAND2_X2 U7972 ( .A1(b[13]), .A2(a[1]), .ZN(n5154) );
  INV_X4 U7973 ( .A(n5154), .ZN(n5156) );
  NAND2_X2 U7974 ( .A1(n5156), .A2(n5155), .ZN(n5196) );
  NAND2_X2 U7975 ( .A1(n5195), .A2(n5196), .ZN(n5158) );
  XNOR2_X2 U7976 ( .A(n5158), .B(n5197), .ZN(n5159) );
  INV_X4 U7977 ( .A(n5159), .ZN(n5306) );
  MUX2_X2 U7978 ( .A(n5161), .B(n5160), .S(n5306), .Z(n5188) );
  XNOR2_X2 U7979 ( .A(n4000), .B(b[14]), .ZN(n5312) );
  XNOR2_X2 U7980 ( .A(n5312), .B(net218392), .ZN(n5311) );
  XNOR2_X2 U7981 ( .A(n5311), .B(net216334), .ZN(n5171) );
  NOR2_X4 U7982 ( .A1(n5162), .A2(n3366), .ZN(n5164) );
  MUX2_X2 U7983 ( .A(net216117), .B(net216517), .S(net218558), .Z(n5163) );
  NAND2_X2 U7984 ( .A1(n5164), .A2(n5163), .ZN(n6982) );
  AOI22_X2 U7985 ( .A1(n7805), .A2(n6278), .B1(n7039), .B2(n6982), .ZN(n5166)
         );
  AOI22_X2 U7986 ( .A1(n7807), .A2(n6272), .B1(n7803), .B2(n5739), .ZN(n5165)
         );
  NAND2_X2 U7987 ( .A1(n5166), .A2(n5165), .ZN(n7811) );
  INV_X4 U7988 ( .A(n7811), .ZN(n5169) );
  NAND2_X2 U7989 ( .A1(n5321), .A2(n5167), .ZN(n5168) );
  AOI21_X2 U7990 ( .B1(n5171), .B2(n3990), .A(n5170), .ZN(n5187) );
  NAND2_X2 U7991 ( .A1(n5327), .A2(n7831), .ZN(n5177) );
  NAND3_X2 U7992 ( .A1(n5177), .A2(n5176), .A3(n5175), .ZN(n5185) );
  INV_X4 U7993 ( .A(n5178), .ZN(n5179) );
  NOR4_X2 U7994 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n5186)
         );
  NAND4_X2 U7995 ( .A1(n5189), .A2(n5188), .A3(n5187), .A4(n5186), .ZN(
        result[14]) );
  NOR2_X4 U7996 ( .A1(n5192), .A2(n5191), .ZN(n5340) );
  NAND2_X2 U7997 ( .A1(n5193), .A2(b[15]), .ZN(n5310) );
  INV_X4 U7998 ( .A(n5195), .ZN(n5198) );
  OAI21_X4 U7999 ( .B1(n5198), .B2(n5197), .A(n5196), .ZN(n5302) );
  INV_X4 U8000 ( .A(n5302), .ZN(n5301) );
  INV_X4 U8001 ( .A(n5199), .ZN(n5203) );
  INV_X4 U8002 ( .A(n5200), .ZN(n5202) );
  OAI21_X4 U8003 ( .B1(n5202), .B2(n5203), .A(n5201), .ZN(n5550) );
  NAND2_X2 U8004 ( .A1(b[13]), .A2(a[2]), .ZN(n5424) );
  XNOR2_X2 U8005 ( .A(n5550), .B(n5424), .ZN(n5299) );
  INV_X4 U8006 ( .A(n5206), .ZN(n5470) );
  INV_X4 U8007 ( .A(n5209), .ZN(n5210) );
  AOI21_X4 U8008 ( .B1(n3416), .B2(n5211), .A(n5210), .ZN(n5469) );
  OAI21_X4 U8009 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n5394) );
  NAND2_X2 U8010 ( .A1(b[8]), .A2(a[7]), .ZN(n5269) );
  INV_X4 U8011 ( .A(n5269), .ZN(n5267) );
  NAND2_X2 U8012 ( .A1(b[7]), .A2(a[8]), .ZN(n5265) );
  INV_X4 U8013 ( .A(n5265), .ZN(n5262) );
  NAND2_X2 U8014 ( .A1(b[6]), .A2(a[9]), .ZN(n5258) );
  INV_X4 U8015 ( .A(n5258), .ZN(n5257) );
  NAND3_X2 U8016 ( .A1(n5219), .A2(net216283), .A3(net216284), .ZN(n5221) );
  INV_X4 U8017 ( .A(n5223), .ZN(n5226) );
  OAI21_X4 U8018 ( .B1(n5226), .B2(n5227), .A(n5225), .ZN(n5356) );
  NAND2_X2 U8019 ( .A1(net218536), .A2(a[12]), .ZN(n5238) );
  INV_X4 U8020 ( .A(n5238), .ZN(n5235) );
  NAND2_X2 U8021 ( .A1(net218548), .A2(a[13]), .ZN(n5228) );
  NAND2_X2 U8022 ( .A1(a[14]), .A2(net218558), .ZN(net216259) );
  NAND2_X2 U8023 ( .A1(n5228), .A2(net216439), .ZN(n5230) );
  INV_X4 U8024 ( .A(net216439), .ZN(net216436) );
  INV_X4 U8025 ( .A(n5228), .ZN(n5229) );
  OAI21_X4 U8026 ( .B1(n5234), .B2(n5233), .A(n5232), .ZN(n5493) );
  XNOR2_X2 U8027 ( .A(n5491), .B(n5493), .ZN(n5236) );
  NAND2_X2 U8028 ( .A1(n5235), .A2(n5236), .ZN(n5367) );
  INV_X4 U8029 ( .A(n5367), .ZN(n5240) );
  INV_X4 U8030 ( .A(n5236), .ZN(n5237) );
  INV_X4 U8031 ( .A(n5364), .ZN(n5239) );
  NOR2_X4 U8032 ( .A1(n5240), .A2(n5239), .ZN(n5248) );
  INV_X4 U8033 ( .A(n5246), .ZN(n5244) );
  XNOR2_X2 U8034 ( .A(n5248), .B(n5247), .ZN(n5249) );
  INV_X4 U8035 ( .A(n5252), .ZN(n5250) );
  NAND2_X2 U8036 ( .A1(b[5]), .A2(a[10]), .ZN(n5251) );
  INV_X4 U8037 ( .A(n5251), .ZN(n5253) );
  NAND2_X2 U8038 ( .A1(n5253), .A2(n5252), .ZN(n5476) );
  NAND2_X2 U8039 ( .A1(n5352), .A2(n5476), .ZN(n5254) );
  XNOR2_X2 U8040 ( .A(n5255), .B(n5254), .ZN(n5259) );
  NAND2_X2 U8041 ( .A1(n5258), .A2(n5259), .ZN(net216220) );
  NAND2_X2 U8042 ( .A1(n5391), .A2(net216220), .ZN(n5260) );
  INV_X4 U8043 ( .A(n5260), .ZN(n5261) );
  XNOR2_X2 U8044 ( .A(n5261), .B(net216400), .ZN(n5263) );
  NAND2_X2 U8045 ( .A1(n5262), .A2(n5263), .ZN(net216022) );
  XNOR2_X2 U8046 ( .A(n5266), .B(net216388), .ZN(n5268) );
  XNOR2_X2 U8047 ( .A(n5272), .B(n5271), .ZN(n5275) );
  INV_X4 U8048 ( .A(n3899), .ZN(n5273) );
  NAND2_X2 U8049 ( .A1(b[9]), .A2(a[6]), .ZN(n5274) );
  INV_X4 U8050 ( .A(n5274), .ZN(n5276) );
  XNOR2_X2 U8051 ( .A(n5278), .B(n5277), .ZN(n5281) );
  INV_X4 U8052 ( .A(n3793), .ZN(n5279) );
  NAND2_X2 U8053 ( .A1(b[10]), .A2(a[5]), .ZN(n5280) );
  INV_X4 U8054 ( .A(n5280), .ZN(n5282) );
  XNOR2_X2 U8055 ( .A(n5284), .B(n5283), .ZN(n5285) );
  NAND2_X2 U8056 ( .A1(b[11]), .A2(net219055), .ZN(n5286) );
  NAND2_X2 U8057 ( .A1(n5285), .A2(n5286), .ZN(n5341) );
  INV_X4 U8058 ( .A(n5286), .ZN(n5542) );
  OAI21_X4 U8059 ( .B1(n5294), .B2(n5293), .A(n5292), .ZN(n5296) );
  XNOR2_X2 U8060 ( .A(n5297), .B(n5342), .ZN(n5551) );
  NAND2_X2 U8061 ( .A1(a[3]), .A2(b[12]), .ZN(n5298) );
  XNOR2_X2 U8062 ( .A(n5299), .B(n5426), .ZN(n5303) );
  NAND2_X2 U8063 ( .A1(n5301), .A2(n5300), .ZN(n5304) );
  NAND2_X2 U8064 ( .A1(n5570), .A2(n5569), .ZN(n5435) );
  INV_X4 U8065 ( .A(n5569), .ZN(n5305) );
  XNOR2_X2 U8066 ( .A(n5307), .B(n5568), .ZN(n5308) );
  INV_X4 U8067 ( .A(n5308), .ZN(n5443) );
  MUX2_X2 U8068 ( .A(n5310), .B(n5309), .S(n5443), .Z(n5339) );
  INV_X4 U8069 ( .A(n5311), .ZN(n5314) );
  INV_X4 U8070 ( .A(n5312), .ZN(n5313) );
  AOI22_X2 U8071 ( .A1(net216334), .A2(n5314), .B1(a[14]), .B2(n5313), .ZN(
        net216128) );
  XNOR2_X2 U8072 ( .A(sel), .B(b[15]), .ZN(net216126) );
  INV_X4 U8073 ( .A(net216129), .ZN(net216332) );
  XNOR2_X2 U8074 ( .A(net216128), .B(net216332), .ZN(n5325) );
  NAND2_X2 U8075 ( .A1(n7803), .A2(n6451), .ZN(n5318) );
  NAND2_X2 U8076 ( .A1(n7807), .A2(n5315), .ZN(n5317) );
  AOI22_X2 U8077 ( .A1(n7039), .A2(net213359), .B1(n7805), .B2(net214477), 
        .ZN(n5316) );
  NAND3_X2 U8078 ( .A1(n5318), .A2(n5317), .A3(n5316), .ZN(n5319) );
  INV_X4 U8079 ( .A(n5319), .ZN(n7876) );
  NAND2_X2 U8080 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  AOI21_X2 U8081 ( .B1(n5325), .B2(n3990), .A(n5324), .ZN(n5338) );
  INV_X4 U8082 ( .A(n7863), .ZN(n5326) );
  NAND2_X2 U8083 ( .A1(n5327), .A2(n5326), .ZN(n5329) );
  NAND3_X2 U8084 ( .A1(n5329), .A2(n7036), .A3(n3409), .ZN(n5336) );
  NOR4_X2 U8085 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n5337)
         );
  NAND4_X2 U8086 ( .A1(n5340), .A2(n5339), .A3(n5338), .A4(n5337), .ZN(
        result[15]) );
  INV_X4 U8087 ( .A(n5342), .ZN(n5343) );
  NAND3_X2 U8088 ( .A1(net216202), .A2(n5396), .A3(n5394), .ZN(net216203) );
  NAND2_X2 U8089 ( .A1(b[7]), .A2(a[9]), .ZN(net216211) );
  INV_X4 U8090 ( .A(net216284), .ZN(net216277) );
  INV_X4 U8091 ( .A(n5359), .ZN(n5366) );
  INV_X4 U8092 ( .A(n5360), .ZN(n5362) );
  NOR3_X4 U8093 ( .A1(n5361), .A2(n5362), .A3(n5366), .ZN(n5369) );
  INV_X4 U8094 ( .A(n5363), .ZN(n5365) );
  OAI21_X4 U8095 ( .B1(n5366), .B2(n5365), .A(n5364), .ZN(n5368) );
  OAI21_X4 U8096 ( .B1(n5369), .B2(n5368), .A(n5367), .ZN(n5485) );
  NAND2_X2 U8097 ( .A1(net218536), .A2(a[13]), .ZN(n5377) );
  INV_X4 U8098 ( .A(net216052), .ZN(net216251) );
  NAND2_X2 U8099 ( .A1(net218548), .A2(a[14]), .ZN(n5495) );
  NAND2_X2 U8100 ( .A1(net216251), .A2(n5495), .ZN(n5494) );
  XNOR2_X2 U8101 ( .A(n5372), .B(n5371), .ZN(n5373) );
  INV_X4 U8102 ( .A(n5377), .ZN(n5374) );
  AOI21_X4 U8103 ( .B1(n5377), .B2(n5376), .A(n5375), .ZN(n5486) );
  XNOR2_X2 U8104 ( .A(n5378), .B(n5486), .ZN(n5381) );
  INV_X4 U8105 ( .A(n5381), .ZN(n5379) );
  NAND2_X2 U8106 ( .A1(b[4]), .A2(a[12]), .ZN(n5380) );
  NAND2_X2 U8107 ( .A1(n5379), .A2(n5380), .ZN(n5482) );
  INV_X4 U8108 ( .A(n5380), .ZN(n5382) );
  NAND2_X2 U8109 ( .A1(n5482), .A2(n5643), .ZN(n5383) );
  XNOR2_X2 U8110 ( .A(n5384), .B(n5383), .ZN(n5385) );
  XNOR2_X2 U8111 ( .A(n5386), .B(n5478), .ZN(n5389) );
  NAND2_X2 U8112 ( .A1(b[6]), .A2(a[10]), .ZN(n5388) );
  INV_X4 U8113 ( .A(n5388), .ZN(n5390) );
  OAI21_X4 U8114 ( .B1(n5392), .B2(net216217), .A(n5391), .ZN(n5475) );
  XNOR2_X2 U8115 ( .A(n5475), .B(n5393), .ZN(net216213) );
  INV_X4 U8116 ( .A(net216213), .ZN(net216212) );
  NAND3_X4 U8117 ( .A1(n5397), .A2(n5396), .A3(net216196), .ZN(net216190) );
  NAND2_X2 U8118 ( .A1(b[9]), .A2(a[7]), .ZN(net216192) );
  INV_X4 U8119 ( .A(net216192), .ZN(net216191) );
  XNOR2_X2 U8120 ( .A(n5399), .B(n5398), .ZN(n5401) );
  NAND2_X2 U8121 ( .A1(b[10]), .A2(a[6]), .ZN(n5400) );
  INV_X4 U8122 ( .A(n5400), .ZN(n5403) );
  XNOR2_X2 U8123 ( .A(n5405), .B(n5404), .ZN(n5408) );
  INV_X4 U8124 ( .A(n5408), .ZN(n5406) );
  NAND2_X2 U8125 ( .A1(b[11]), .A2(a[5]), .ZN(n5407) );
  INV_X4 U8126 ( .A(n5407), .ZN(n5409) );
  XNOR2_X2 U8127 ( .A(n5411), .B(n5410), .ZN(n5414) );
  NAND2_X2 U8128 ( .A1(b[12]), .A2(net219055), .ZN(n5413) );
  INV_X4 U8129 ( .A(n5413), .ZN(n5415) );
  INV_X4 U8130 ( .A(n5624), .ZN(n5417) );
  XNOR2_X2 U8131 ( .A(n5419), .B(n5418), .ZN(n5422) );
  NAND2_X2 U8132 ( .A1(b[13]), .A2(a[3]), .ZN(n5421) );
  INV_X4 U8133 ( .A(n5421), .ZN(n5423) );
  INV_X4 U8134 ( .A(n5424), .ZN(n5428) );
  NAND2_X2 U8135 ( .A1(n5425), .A2(n5624), .ZN(n5426) );
  NAND2_X2 U8136 ( .A1(n5428), .A2(n5427), .ZN(n5616) );
  XNOR2_X2 U8137 ( .A(n5430), .B(n5429), .ZN(n5433) );
  NAND2_X2 U8138 ( .A1(b[14]), .A2(a[2]), .ZN(n5432) );
  INV_X4 U8139 ( .A(n5432), .ZN(n5434) );
  NAND2_X2 U8140 ( .A1(n5434), .A2(n5433), .ZN(n5575) );
  NAND2_X2 U8141 ( .A1(n5574), .A2(n5575), .ZN(n5438) );
  INV_X4 U8142 ( .A(n5435), .ZN(n5436) );
  XNOR2_X2 U8143 ( .A(n5438), .B(n5437), .ZN(n5441) );
  INV_X4 U8144 ( .A(n5441), .ZN(n5439) );
  INV_X4 U8145 ( .A(n5440), .ZN(n5442) );
  NAND3_X4 U8146 ( .A1(a[0]), .A2(b[15]), .A3(n5443), .ZN(n5582) );
  XNOR2_X2 U8147 ( .A(n5444), .B(n5582), .ZN(n5445) );
  INV_X4 U8148 ( .A(n5445), .ZN(n5588) );
  OAI211_X2 U8149 ( .C1(n5588), .C2(n7888), .A(net218608), .B(n3400), .ZN(
        n5448) );
  NAND2_X2 U8150 ( .A1(n5446), .A2(n7807), .ZN(n6983) );
  AOI21_X2 U8151 ( .B1(b[16]), .B2(n5448), .A(n5447), .ZN(n5468) );
  NAND2_X2 U8152 ( .A1(n7033), .A2(n5449), .ZN(n5467) );
  INV_X4 U8153 ( .A(b[16]), .ZN(net216135) );
  NAND2_X2 U8154 ( .A1(net218658), .A2(net216135), .ZN(n5450) );
  NAND2_X2 U8155 ( .A1(n5450), .A2(net212094), .ZN(n5452) );
  NAND2_X2 U8156 ( .A1(n7821), .A2(b[4]), .ZN(n7058) );
  INV_X4 U8157 ( .A(n7058), .ZN(n6101) );
  NAND2_X2 U8158 ( .A1(n6101), .A2(n7039), .ZN(n6454) );
  INV_X4 U8159 ( .A(n6454), .ZN(n5736) );
  XNOR2_X2 U8160 ( .A(n4000), .B(b[16]), .ZN(n5599) );
  XNOR2_X2 U8161 ( .A(n5599), .B(net216124), .ZN(n5598) );
  XNOR2_X2 U8162 ( .A(n5598), .B(net215913), .ZN(n5464) );
  NAND2_X2 U8163 ( .A1(net218639), .A2(n5453), .ZN(n5454) );
  OAI211_X2 U8164 ( .C1(n6653), .C2(n5455), .A(n5454), .B(n3401), .ZN(n5463)
         );
  MUX2_X2 U8165 ( .A(net215701), .B(net216117), .S(net218556), .Z(n5457) );
  NAND2_X2 U8166 ( .A1(n5458), .A2(n5457), .ZN(n6630) );
  NAND2_X2 U8167 ( .A1(n7050), .A2(n6630), .ZN(n5461) );
  NAND2_X2 U8168 ( .A1(n6851), .A2(n5459), .ZN(n5460) );
  NAND2_X2 U8169 ( .A1(n5461), .A2(n5460), .ZN(n5462) );
  AOI211_X2 U8170 ( .C1(n5464), .C2(n3990), .A(n5463), .B(n5462), .ZN(n5465)
         );
  NAND4_X2 U8171 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(
        result[16]) );
  NAND2_X2 U8172 ( .A1(a[3]), .A2(b[14]), .ZN(n5566) );
  INV_X4 U8173 ( .A(n5566), .ZN(n5564) );
  NAND2_X2 U8174 ( .A1(b[13]), .A2(net219055), .ZN(n5559) );
  INV_X4 U8175 ( .A(n5559), .ZN(n5557) );
  NAND2_X2 U8176 ( .A1(b[12]), .A2(a[5]), .ZN(n5548) );
  INV_X4 U8177 ( .A(n5548), .ZN(n5547) );
  NAND2_X2 U8178 ( .A1(b[10]), .A2(a[7]), .ZN(n5529) );
  INV_X4 U8179 ( .A(n5529), .ZN(n5527) );
  OAI21_X4 U8180 ( .B1(n3980), .B2(n5478), .A(n3175), .ZN(n5479) );
  INV_X4 U8181 ( .A(n5480), .ZN(n5484) );
  INV_X4 U8182 ( .A(n5481), .ZN(n5483) );
  OAI21_X4 U8183 ( .B1(n5483), .B2(n5484), .A(n5482), .ZN(n5644) );
  NAND2_X2 U8184 ( .A1(net218536), .A2(a[14]), .ZN(n5503) );
  NAND2_X2 U8185 ( .A1(net218548), .A2(a[15]), .ZN(n5487) );
  NAND2_X2 U8186 ( .A1(net216064), .A2(n5487), .ZN(n5654) );
  INV_X4 U8187 ( .A(n5487), .ZN(n5488) );
  INV_X4 U8188 ( .A(net216064), .ZN(net216063) );
  NAND2_X2 U8189 ( .A1(n5654), .A2(n5783), .ZN(n5501) );
  INV_X4 U8190 ( .A(n5495), .ZN(n5490) );
  INV_X4 U8191 ( .A(n5496), .ZN(n5489) );
  NAND2_X2 U8192 ( .A1(n5490), .A2(n5489), .ZN(n5500) );
  INV_X4 U8193 ( .A(n5491), .ZN(n5492) );
  NAND3_X2 U8194 ( .A1(n5494), .A2(n5493), .A3(n5492), .ZN(n5499) );
  NAND2_X2 U8195 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  NAND2_X2 U8196 ( .A1(net216052), .A2(n5497), .ZN(n5498) );
  NAND3_X2 U8197 ( .A1(n5500), .A2(n5499), .A3(n5498), .ZN(n5655) );
  XNOR2_X2 U8198 ( .A(n5501), .B(n5655), .ZN(n5504) );
  NAND2_X2 U8199 ( .A1(n5503), .A2(n5502), .ZN(n5505) );
  NAND3_X2 U8200 ( .A1(a[14]), .A2(n5504), .A3(net218536), .ZN(n5779) );
  XNOR2_X2 U8201 ( .A(n5506), .B(n5651), .ZN(n5507) );
  XNOR2_X2 U8202 ( .A(n5508), .B(n5645), .ZN(n5509) );
  XNOR2_X2 U8203 ( .A(n5805), .B(n5510), .ZN(n5513) );
  NAND2_X2 U8204 ( .A1(b[6]), .A2(a[11]), .ZN(n5512) );
  INV_X4 U8205 ( .A(n5512), .ZN(n5514) );
  NAND2_X2 U8206 ( .A1(b[7]), .A2(a[10]), .ZN(n5517) );
  INV_X4 U8207 ( .A(n5517), .ZN(n5518) );
  NAND2_X2 U8208 ( .A1(n5518), .A2(n3946), .ZN(net215814) );
  NAND2_X2 U8209 ( .A1(b[9]), .A2(a[8]), .ZN(n5519) );
  INV_X4 U8210 ( .A(n5519), .ZN(n5520) );
  XNOR2_X2 U8211 ( .A(n5526), .B(n5688), .ZN(n5528) );
  INV_X4 U8212 ( .A(n5528), .ZN(n5530) );
  XNOR2_X2 U8213 ( .A(n5532), .B(n5531), .ZN(n5535) );
  NAND2_X2 U8214 ( .A1(b[11]), .A2(a[6]), .ZN(n5534) );
  INV_X4 U8215 ( .A(n5534), .ZN(n5536) );
  INV_X4 U8216 ( .A(n5537), .ZN(n5546) );
  NAND2_X2 U8217 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  AOI21_X4 U8218 ( .B1(n5544), .B2(n5633), .A(n5543), .ZN(n5545) );
  INV_X4 U8219 ( .A(n5549), .ZN(n5556) );
  XNOR2_X2 U8220 ( .A(n5556), .B(n5555), .ZN(n5558) );
  NAND2_X2 U8221 ( .A1(b[15]), .A2(a[2]), .ZN(n5716) );
  XNOR2_X2 U8222 ( .A(n5567), .B(n5716), .ZN(n5578) );
  NOR2_X4 U8223 ( .A1(n5573), .A2(n5572), .ZN(n5577) );
  INV_X4 U8224 ( .A(n5574), .ZN(n5576) );
  OAI21_X4 U8225 ( .B1(n5576), .B2(n5577), .A(n5575), .ZN(n5846) );
  XNOR2_X2 U8226 ( .A(n5578), .B(n3932), .ZN(n5889) );
  INV_X4 U8227 ( .A(n5582), .ZN(n5579) );
  INV_X4 U8228 ( .A(n5580), .ZN(n5769) );
  INV_X4 U8229 ( .A(n5581), .ZN(n5583) );
  OAI21_X4 U8230 ( .B1(n5583), .B2(n5582), .A(net215476), .ZN(n5715) );
  NAND2_X2 U8231 ( .A1(b[16]), .A2(a[1]), .ZN(n5584) );
  INV_X4 U8232 ( .A(n5584), .ZN(n5587) );
  NAND3_X4 U8233 ( .A1(a[0]), .A2(b[16]), .A3(n5588), .ZN(n5761) );
  XNOR2_X2 U8234 ( .A(n5589), .B(n5761), .ZN(n5592) );
  INV_X4 U8235 ( .A(n5592), .ZN(n5732) );
  OAI211_X2 U8236 ( .C1(n5732), .C2(net218655), .A(net218608), .B(n3412), .ZN(
        n5594) );
  AOI211_X4 U8237 ( .C1(b[17]), .C2(n5594), .A(n5593), .B(n3384), .ZN(n5613)
         );
  INV_X4 U8238 ( .A(n6983), .ZN(n7031) );
  NAND4_X2 U8239 ( .A1(n5597), .A2(net215919), .A3(net215920), .A4(n5596), 
        .ZN(n6849) );
  INV_X4 U8240 ( .A(n6849), .ZN(n7221) );
  INV_X4 U8241 ( .A(n5598), .ZN(n5601) );
  INV_X4 U8242 ( .A(n5599), .ZN(n5600) );
  AOI22_X2 U8243 ( .A1(net215913), .A2(n5601), .B1(a[16]), .B2(n5600), .ZN(
        n5741) );
  XNOR2_X2 U8244 ( .A(sel), .B(b[17]), .ZN(n5742) );
  XNOR2_X2 U8245 ( .A(n5742), .B(net218378), .ZN(n5740) );
  XNOR2_X2 U8246 ( .A(n5741), .B(n5740), .ZN(n5604) );
  INV_X4 U8247 ( .A(n7035), .ZN(n6468) );
  NAND2_X2 U8248 ( .A1(n6468), .A2(n5602), .ZN(n5603) );
  OAI221_X2 U8249 ( .B1(n7221), .B2(n6135), .C1(n7389), .C2(n5604), .A(n5603), 
        .ZN(n5610) );
  NAND2_X2 U8250 ( .A1(net218639), .A2(n5605), .ZN(n5606) );
  NOR3_X2 U8251 ( .A1(n5610), .A2(n5609), .A3(n5608), .ZN(n5611) );
  NAND3_X2 U8252 ( .A1(n5613), .A2(n5612), .A3(n5611), .ZN(result[17]) );
  NAND2_X2 U8253 ( .A1(b[17]), .A2(a[1]), .ZN(n5730) );
  INV_X4 U8254 ( .A(n5634), .ZN(n5635) );
  NAND2_X2 U8255 ( .A1(b[7]), .A2(a[11]), .ZN(n5684) );
  INV_X4 U8256 ( .A(n5684), .ZN(n5682) );
  OAI21_X4 U8257 ( .B1(n5642), .B2(n5641), .A(n5640), .ZN(n5771) );
  INV_X4 U8258 ( .A(n5643), .ZN(n5648) );
  INV_X4 U8259 ( .A(n5644), .ZN(n5647) );
  OAI21_X4 U8260 ( .B1(n5647), .B2(n5648), .A(n5646), .ZN(n5799) );
  INV_X4 U8261 ( .A(n5650), .ZN(n5653) );
  INV_X4 U8262 ( .A(n5651), .ZN(n5652) );
  OAI21_X4 U8263 ( .B1(n5375), .B2(n5653), .A(n5652), .ZN(n5778) );
  NAND2_X2 U8264 ( .A1(n5778), .A2(n5779), .ZN(n5663) );
  NAND2_X2 U8265 ( .A1(net218536), .A2(a[15]), .ZN(n5660) );
  NAND2_X2 U8266 ( .A1(net218548), .A2(a[16]), .ZN(n5656) );
  INV_X4 U8267 ( .A(net215846), .ZN(net215848) );
  NAND3_X2 U8268 ( .A1(a[16]), .A2(net215846), .A3(net218548), .ZN(n5920) );
  NAND2_X2 U8269 ( .A1(n5785), .A2(n5920), .ZN(n5657) );
  XNOR2_X2 U8270 ( .A(n5658), .B(n5657), .ZN(n5661) );
  INV_X4 U8271 ( .A(n5661), .ZN(n5659) );
  XNOR2_X2 U8272 ( .A(n5663), .B(n5777), .ZN(n5666) );
  INV_X4 U8273 ( .A(n5666), .ZN(n5664) );
  NAND2_X2 U8274 ( .A1(a[14]), .A2(b[4]), .ZN(n5665) );
  INV_X4 U8275 ( .A(n5665), .ZN(n5667) );
  NAND2_X2 U8276 ( .A1(n5667), .A2(n3908), .ZN(n5795) );
  NAND2_X2 U8277 ( .A1(n5796), .A2(n5795), .ZN(n5668) );
  XNOR2_X2 U8278 ( .A(n5669), .B(n5668), .ZN(n5672) );
  INV_X4 U8279 ( .A(n5672), .ZN(n5670) );
  NAND2_X2 U8280 ( .A1(a[13]), .A2(b[5]), .ZN(n5671) );
  INV_X4 U8281 ( .A(n5671), .ZN(n5673) );
  XNOR2_X2 U8282 ( .A(n5947), .B(n5674), .ZN(n5678) );
  INV_X4 U8283 ( .A(n5678), .ZN(n5676) );
  NAND2_X2 U8284 ( .A1(b[6]), .A2(a[12]), .ZN(n5677) );
  INV_X4 U8285 ( .A(n5677), .ZN(n5679) );
  XNOR2_X2 U8286 ( .A(n5681), .B(n5680), .ZN(n5683) );
  XNOR2_X2 U8287 ( .A(net219656), .B(net215805), .ZN(n5687) );
  INV_X4 U8288 ( .A(n5687), .ZN(n5686) );
  NAND2_X2 U8289 ( .A1(b[8]), .A2(a[10]), .ZN(net215802) );
  INV_X4 U8290 ( .A(net215777), .ZN(net215781) );
  NAND2_X2 U8291 ( .A1(b[10]), .A2(a[8]), .ZN(n5689) );
  OAI21_X4 U8292 ( .B1(net215780), .B2(net215781), .A(n5689), .ZN(n5911) );
  INV_X4 U8293 ( .A(n5689), .ZN(n5690) );
  XNOR2_X2 U8294 ( .A(net215775), .B(net215776), .ZN(n5692) );
  NAND2_X2 U8295 ( .A1(b[11]), .A2(a[7]), .ZN(net215773) );
  XNOR2_X2 U8296 ( .A(n5693), .B(net215770), .ZN(n5696) );
  INV_X4 U8297 ( .A(n5696), .ZN(n5694) );
  NAND2_X2 U8298 ( .A1(b[12]), .A2(a[6]), .ZN(n5695) );
  INV_X4 U8299 ( .A(n5695), .ZN(n5697) );
  XNOR2_X2 U8300 ( .A(n5699), .B(n5698), .ZN(n5702) );
  INV_X4 U8301 ( .A(n5702), .ZN(n5700) );
  NAND2_X2 U8302 ( .A1(b[13]), .A2(a[5]), .ZN(n5701) );
  INV_X4 U8303 ( .A(n5701), .ZN(n5703) );
  XNOR2_X2 U8304 ( .A(n5705), .B(n5704), .ZN(n5707) );
  NAND2_X2 U8305 ( .A1(b[14]), .A2(net219055), .ZN(n5706) );
  INV_X4 U8306 ( .A(n5706), .ZN(n5708) );
  XNOR2_X2 U8307 ( .A(n5710), .B(n5709), .ZN(n5713) );
  NAND2_X2 U8308 ( .A1(a[3]), .A2(b[15]), .ZN(n5712) );
  INV_X4 U8309 ( .A(n5712), .ZN(n5714) );
  NAND2_X2 U8310 ( .A1(n5714), .A2(n5713), .ZN(net215471) );
  INV_X4 U8311 ( .A(n5715), .ZN(n5720) );
  INV_X4 U8312 ( .A(n5716), .ZN(n5719) );
  XNOR2_X2 U8313 ( .A(n5722), .B(n5721), .ZN(n5724) );
  NAND2_X2 U8314 ( .A1(b[16]), .A2(a[2]), .ZN(n5723) );
  INV_X4 U8315 ( .A(n5723), .ZN(n5725) );
  NAND2_X2 U8316 ( .A1(n5760), .A2(n5766), .ZN(n5728) );
  INV_X4 U8317 ( .A(n5764), .ZN(n5726) );
  XNOR2_X2 U8318 ( .A(n5728), .B(n5727), .ZN(n5731) );
  INV_X4 U8319 ( .A(n5731), .ZN(n5729) );
  NAND3_X4 U8320 ( .A1(a[0]), .A2(b[17]), .A3(n5732), .ZN(n5757) );
  NOR2_X4 U8321 ( .A1(net212677), .A2(n5733), .ZN(n5734) );
  OAI21_X4 U8322 ( .B1(n5735), .B2(n5734), .A(n7036), .ZN(n5737) );
  AOI211_X4 U8323 ( .C1(b[18]), .C2(n5738), .A(n5737), .B(n3382), .ZN(n5756)
         );
  XNOR2_X2 U8324 ( .A(n4002), .B(b[18]), .ZN(n5871) );
  OAI22_X2 U8325 ( .A1(n5742), .A2(net218378), .B1(n5741), .B2(n5740), .ZN(
        n5873) );
  XNOR2_X2 U8326 ( .A(n3334), .B(n5873), .ZN(n5744) );
  NAND2_X2 U8327 ( .A1(net218639), .A2(n3378), .ZN(n5743) );
  OAI211_X2 U8328 ( .C1(n7389), .C2(n5744), .A(n5743), .B(n3399), .ZN(n5753)
         );
  INV_X4 U8329 ( .A(n5745), .ZN(n5751) );
  NOR2_X4 U8330 ( .A1(n5746), .A2(n3367), .ZN(n5748) );
  MUX2_X2 U8331 ( .A(net215245), .B(net215701), .S(net218556), .Z(n5747) );
  NAND2_X2 U8332 ( .A1(n5748), .A2(n5747), .ZN(n7806) );
  NAND2_X2 U8333 ( .A1(n7050), .A2(n7806), .ZN(n5749) );
  OAI221_X2 U8334 ( .B1(n5751), .B2(n7035), .C1(n5750), .C2(n6637), .A(n5749), 
        .ZN(n5752) );
  NOR2_X2 U8335 ( .A1(n5753), .A2(n5752), .ZN(n5754) );
  NAND3_X2 U8336 ( .A1(n5756), .A2(n5755), .A3(n5754), .ZN(result[18]) );
  INV_X4 U8337 ( .A(n5757), .ZN(n5759) );
  INV_X4 U8338 ( .A(n5863), .ZN(n5858) );
  INV_X4 U8339 ( .A(n5760), .ZN(n5768) );
  INV_X4 U8340 ( .A(n5761), .ZN(n5765) );
  INV_X4 U8341 ( .A(n5762), .ZN(n5763) );
  AOI21_X4 U8342 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(n5767) );
  OAI21_X4 U8343 ( .B1(n5768), .B2(n5767), .A(n5766), .ZN(n6012) );
  NAND2_X2 U8344 ( .A1(b[15]), .A2(net219055), .ZN(n5852) );
  INV_X4 U8345 ( .A(n5852), .ZN(n5851) );
  NAND2_X2 U8346 ( .A1(b[14]), .A2(a[5]), .ZN(n5842) );
  INV_X4 U8347 ( .A(n5842), .ZN(n5840) );
  NAND2_X2 U8348 ( .A1(b[13]), .A2(a[6]), .ZN(n5835) );
  NAND2_X2 U8349 ( .A1(b[12]), .A2(a[7]), .ZN(n5826) );
  INV_X4 U8350 ( .A(n5826), .ZN(n5824) );
  NAND2_X2 U8351 ( .A1(b[11]), .A2(a[8]), .ZN(net215568) );
  NAND2_X2 U8352 ( .A1(b[10]), .A2(a[9]), .ZN(n5821) );
  INV_X4 U8353 ( .A(n5821), .ZN(n5819) );
  NAND2_X2 U8354 ( .A1(n3605), .A2(n5771), .ZN(n5775) );
  AOI21_X4 U8355 ( .B1(n5776), .B2(n5775), .A(n5774), .ZN(n5958) );
  AOI21_X4 U8356 ( .B1(n5779), .B2(n5778), .A(n5777), .ZN(n5782) );
  INV_X4 U8357 ( .A(n5780), .ZN(n5781) );
  NOR2_X4 U8358 ( .A1(n5782), .A2(n5781), .ZN(n5934) );
  NAND2_X2 U8359 ( .A1(net218536), .A2(a[16]), .ZN(n5790) );
  NAND2_X2 U8360 ( .A1(n5658), .A2(n5785), .ZN(n5921) );
  NAND2_X2 U8361 ( .A1(net218548), .A2(a[17]), .ZN(n5786) );
  NAND2_X2 U8362 ( .A1(a[18]), .A2(net218558), .ZN(net215424) );
  NAND2_X2 U8363 ( .A1(n5786), .A2(net215636), .ZN(n5922) );
  INV_X4 U8364 ( .A(net215636), .ZN(net215635) );
  NAND2_X2 U8365 ( .A1(n5922), .A2(n5919), .ZN(n5787) );
  XNOR2_X2 U8366 ( .A(n5788), .B(n5787), .ZN(n5791) );
  INV_X4 U8367 ( .A(n5791), .ZN(n5789) );
  NAND2_X2 U8368 ( .A1(n5790), .A2(n5789), .ZN(n5792) );
  NAND3_X2 U8369 ( .A1(a[16]), .A2(n5791), .A3(net218536), .ZN(n5932) );
  NAND2_X2 U8370 ( .A1(n5792), .A2(n5932), .ZN(n5933) );
  INV_X4 U8371 ( .A(n5933), .ZN(n5793) );
  XNOR2_X2 U8372 ( .A(n5934), .B(n5793), .ZN(n5794) );
  INV_X4 U8373 ( .A(n5795), .ZN(n5937) );
  INV_X4 U8374 ( .A(n5796), .ZN(n5797) );
  AOI21_X4 U8375 ( .B1(n5799), .B2(n5798), .A(n5797), .ZN(n5936) );
  NOR2_X4 U8376 ( .A1(n5936), .A2(n5937), .ZN(n5800) );
  XNOR2_X2 U8377 ( .A(n5801), .B(n5800), .ZN(n5946) );
  NAND2_X2 U8378 ( .A1(a[14]), .A2(b[5]), .ZN(n5942) );
  INV_X4 U8379 ( .A(n5948), .ZN(n5807) );
  OAI21_X4 U8380 ( .B1(n5805), .B2(n3786), .A(n3572), .ZN(n5947) );
  INV_X4 U8381 ( .A(n5947), .ZN(n5806) );
  OAI21_X4 U8382 ( .B1(n5806), .B2(n5807), .A(n3930), .ZN(n5808) );
  XNOR2_X2 U8383 ( .A(n5809), .B(n5808), .ZN(n5810) );
  XNOR2_X2 U8384 ( .A(n5958), .B(n5811), .ZN(n5814) );
  NAND2_X2 U8385 ( .A1(b[7]), .A2(a[12]), .ZN(n5813) );
  INV_X4 U8386 ( .A(n5813), .ZN(n5815) );
  XNOR2_X2 U8387 ( .A(n5817), .B(n5816), .ZN(net215431) );
  NAND2_X2 U8388 ( .A1(b[8]), .A2(a[11]), .ZN(net215595) );
  XNOR2_X2 U8389 ( .A(n5818), .B(net215593), .ZN(net215589) );
  INV_X4 U8390 ( .A(net215589), .ZN(net215591) );
  NAND2_X2 U8391 ( .A1(b[9]), .A2(a[10]), .ZN(net215590) );
  XNOR2_X2 U8392 ( .A(net215581), .B(net215582), .ZN(n5820) );
  XNOR2_X2 U8393 ( .A(net215571), .B(n5823), .ZN(net215569) );
  XNOR2_X2 U8394 ( .A(net215566), .B(net215565), .ZN(n5825) );
  NAND2_X2 U8395 ( .A1(n5824), .A2(n5825), .ZN(n6020) );
  NAND2_X2 U8396 ( .A1(n5906), .A2(n6020), .ZN(n5828) );
  INV_X4 U8397 ( .A(n5828), .ZN(n5832) );
  AOI21_X4 U8398 ( .B1(n5830), .B2(n5907), .A(n5829), .ZN(n5831) );
  XNOR2_X2 U8399 ( .A(n5832), .B(n5831), .ZN(n5834) );
  INV_X4 U8400 ( .A(n5901), .ZN(n6019) );
  INV_X4 U8401 ( .A(n3906), .ZN(n5836) );
  NOR2_X4 U8402 ( .A1(n6019), .A2(n5836), .ZN(n5839) );
  INV_X4 U8403 ( .A(n5897), .ZN(n5837) );
  AOI21_X2 U8404 ( .B1(n5705), .B2(n5900), .A(n5837), .ZN(n5838) );
  INV_X4 U8405 ( .A(n5844), .ZN(n5850) );
  XNOR2_X2 U8406 ( .A(n5853), .B(net215530), .ZN(n5854) );
  INV_X4 U8407 ( .A(n6013), .ZN(n5855) );
  NAND2_X2 U8408 ( .A1(a[3]), .A2(b[16]), .ZN(n5856) );
  INV_X4 U8409 ( .A(n5856), .ZN(n6014) );
  XNOR2_X2 U8410 ( .A(n5857), .B(n5973), .ZN(n5860) );
  OAI21_X4 U8411 ( .B1(n5859), .B2(n5858), .A(n5860), .ZN(net214732) );
  INV_X4 U8412 ( .A(net215516), .ZN(net215519) );
  NAND2_X2 U8413 ( .A1(b[18]), .A2(a[1]), .ZN(net215518) );
  INV_X4 U8414 ( .A(net215518), .ZN(net215517) );
  NAND2_X2 U8415 ( .A1(net215282), .A2(n5980), .ZN(n5864) );
  INV_X4 U8416 ( .A(n5867), .ZN(n5984) );
  OAI211_X2 U8417 ( .C1(n5984), .C2(n7888), .A(net218608), .B(n3403), .ZN(
        n5870) );
  AOI211_X4 U8418 ( .C1(b[19]), .C2(n5870), .A(n5869), .B(n5868), .ZN(n5885)
         );
  INV_X4 U8419 ( .A(n5871), .ZN(n5872) );
  AOI22_X2 U8420 ( .A1(n5873), .A2(n3334), .B1(a[18]), .B2(n5872), .ZN(n5996)
         );
  XNOR2_X2 U8421 ( .A(sel), .B(b[19]), .ZN(n5997) );
  XNOR2_X2 U8422 ( .A(n5997), .B(net215499), .ZN(n5995) );
  XNOR2_X2 U8423 ( .A(n5996), .B(n5995), .ZN(n5876) );
  NAND2_X2 U8424 ( .A1(net218639), .A2(n5874), .ZN(n5875) );
  OAI211_X2 U8425 ( .C1(n7389), .C2(n5876), .A(n5875), .B(n3404), .ZN(n5882)
         );
  NAND2_X2 U8426 ( .A1(n7050), .A2(net212010), .ZN(n5879) );
  INV_X4 U8427 ( .A(n6637), .ZN(n7040) );
  NAND2_X2 U8428 ( .A1(n7040), .A2(n5877), .ZN(n5878) );
  OAI211_X2 U8429 ( .C1(n5880), .C2(n7035), .A(n5879), .B(n5878), .ZN(n5881)
         );
  NOR2_X2 U8430 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  NAND3_X2 U8431 ( .A1(n5885), .A2(n5884), .A3(n5883), .ZN(result[19]) );
  NAND2_X2 U8432 ( .A1(a[3]), .A2(b[17]), .ZN(net215294) );
  INV_X4 U8433 ( .A(net215294), .ZN(net215296) );
  INV_X4 U8434 ( .A(n5886), .ZN(n5887) );
  NAND3_X2 U8435 ( .A1(n5896), .A2(n5897), .A3(n5898), .ZN(n5899) );
  NAND3_X4 U8436 ( .A1(n5900), .A2(n3906), .A3(n5899), .ZN(n6017) );
  NAND3_X2 U8437 ( .A1(n5907), .A2(n5906), .A3(n5905), .ZN(n6021) );
  OAI21_X4 U8438 ( .B1(n5916), .B2(n3787), .A(net215434), .ZN(net215334) );
  NAND2_X2 U8439 ( .A1(net218536), .A2(a[17]), .ZN(n5929) );
  NAND2_X2 U8440 ( .A1(net218548), .A2(a[18]), .ZN(n5917) );
  INV_X4 U8441 ( .A(net215414), .ZN(net215416) );
  NAND2_X2 U8442 ( .A1(n5917), .A2(net215416), .ZN(n5918) );
  NAND3_X2 U8443 ( .A1(a[18]), .A2(net215414), .A3(net218548), .ZN(n6035) );
  INV_X4 U8444 ( .A(n6036), .ZN(n5927) );
  INV_X4 U8445 ( .A(n5919), .ZN(n6034) );
  INV_X4 U8446 ( .A(n5921), .ZN(n5923) );
  OAI21_X4 U8447 ( .B1(n5924), .B2(n5923), .A(n5922), .ZN(n5925) );
  INV_X4 U8448 ( .A(n5925), .ZN(n6033) );
  NOR2_X4 U8449 ( .A1(n6034), .A2(n6033), .ZN(n5926) );
  XNOR2_X2 U8450 ( .A(n5927), .B(n5926), .ZN(n5930) );
  NAND2_X2 U8451 ( .A1(n5929), .A2(n5928), .ZN(n5931) );
  NAND3_X2 U8452 ( .A1(a[17]), .A2(n5930), .A3(net218536), .ZN(n6044) );
  OAI21_X4 U8453 ( .B1(n5934), .B2(n5933), .A(n5932), .ZN(n6043) );
  XNOR2_X2 U8454 ( .A(n6045), .B(n6043), .ZN(n5935) );
  OAI21_X4 U8455 ( .B1(n3310), .B2(n3788), .A(n6050), .ZN(n6051) );
  NOR2_X4 U8456 ( .A1(n5937), .A2(n5936), .ZN(n5940) );
  XNOR2_X2 U8457 ( .A(n6051), .B(n6049), .ZN(n5941) );
  NAND2_X2 U8458 ( .A1(n5943), .A2(n5942), .ZN(n5945) );
  NAND2_X2 U8459 ( .A1(n5951), .A2(n5950), .ZN(n6031) );
  XNOR2_X2 U8460 ( .A(n6030), .B(n6031), .ZN(n5954) );
  INV_X4 U8461 ( .A(n5954), .ZN(n5952) );
  NAND2_X2 U8462 ( .A1(a[14]), .A2(b[6]), .ZN(n5953) );
  NAND2_X2 U8463 ( .A1(n5952), .A2(n5953), .ZN(n6029) );
  INV_X4 U8464 ( .A(n5953), .ZN(n5955) );
  NAND2_X2 U8465 ( .A1(n5955), .A2(n5954), .ZN(n6157) );
  NAND2_X2 U8466 ( .A1(n6029), .A2(n6157), .ZN(n5960) );
  XNOR2_X2 U8467 ( .A(n5960), .B(n5959), .ZN(n6024) );
  NAND2_X2 U8468 ( .A1(b[7]), .A2(a[13]), .ZN(net215206) );
  AOI21_X4 U8469 ( .B1(n5817), .B2(n6026), .A(n6022), .ZN(net215360) );
  NAND2_X2 U8470 ( .A1(b[8]), .A2(a[12]), .ZN(net215357) );
  XNOR2_X2 U8471 ( .A(net215327), .B(net215328), .ZN(net215324) );
  NAND2_X2 U8472 ( .A1(b[12]), .A2(a[8]), .ZN(net215325) );
  NAND2_X2 U8473 ( .A1(b[13]), .A2(a[7]), .ZN(n5963) );
  INV_X4 U8474 ( .A(n5963), .ZN(n5964) );
  NAND2_X2 U8475 ( .A1(n5964), .A2(net215318), .ZN(net214971) );
  XNOR2_X2 U8476 ( .A(n5965), .B(net215316), .ZN(n5968) );
  INV_X4 U8477 ( .A(n5968), .ZN(n5966) );
  NAND2_X2 U8478 ( .A1(b[14]), .A2(a[6]), .ZN(n5967) );
  INV_X4 U8479 ( .A(n5967), .ZN(n5969) );
  NAND2_X2 U8480 ( .A1(n3883), .A2(n5969), .ZN(net215090) );
  NAND2_X2 U8481 ( .A1(b[15]), .A2(a[5]), .ZN(net215307) );
  XNOR2_X2 U8482 ( .A(n5970), .B(net215298), .ZN(net215295) );
  INV_X4 U8483 ( .A(n3920), .ZN(n5971) );
  INV_X4 U8484 ( .A(n5972), .ZN(n5975) );
  XNOR2_X2 U8485 ( .A(net215287), .B(n6300), .ZN(n5978) );
  NAND2_X2 U8486 ( .A1(b[18]), .A2(a[2]), .ZN(n5977) );
  INV_X4 U8487 ( .A(n5977), .ZN(n5979) );
  INV_X4 U8488 ( .A(net215282), .ZN(net215279) );
  OAI21_X4 U8489 ( .B1(net215279), .B2(n5981), .A(n5980), .ZN(net215058) );
  INV_X4 U8490 ( .A(net215275), .ZN(net215277) );
  NAND2_X2 U8491 ( .A1(b[19]), .A2(a[1]), .ZN(n5982) );
  INV_X4 U8492 ( .A(n5982), .ZN(n5983) );
  NAND3_X4 U8493 ( .A1(a[0]), .A2(b[19]), .A3(n5984), .ZN(n6088) );
  XNOR2_X2 U8494 ( .A(n5985), .B(n6088), .ZN(n5988) );
  INV_X4 U8495 ( .A(n5988), .ZN(n6097) );
  INV_X4 U8496 ( .A(n6630), .ZN(n7074) );
  NOR3_X4 U8497 ( .A1(n5994), .A2(n5993), .A3(n5992), .ZN(n6010) );
  XNOR2_X2 U8498 ( .A(n4002), .B(b[20]), .ZN(n6105) );
  INV_X4 U8499 ( .A(a[19]), .ZN(net215256) );
  OAI22_X2 U8500 ( .A1(n5997), .A2(net215256), .B1(n5996), .B2(n5995), .ZN(
        n6107) );
  XNOR2_X2 U8501 ( .A(n3335), .B(n6107), .ZN(n6000) );
  NAND2_X2 U8502 ( .A1(net218639), .A2(n5998), .ZN(n5999) );
  OAI211_X2 U8503 ( .C1(n7389), .C2(n6000), .A(n5999), .B(n3402), .ZN(n6008)
         );
  MUX2_X2 U8504 ( .A(net215001), .B(net215245), .S(net218558), .Z(n6002) );
  NOR2_X2 U8505 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  NAND2_X2 U8506 ( .A1(net218658), .A2(net215232), .ZN(n6099) );
  OAI21_X4 U8507 ( .B1(n5888), .B2(n6016), .A(n6015), .ZN(net214720) );
  NAND2_X2 U8508 ( .A1(n6021), .A2(n6020), .ZN(net215218) );
  NAND2_X2 U8509 ( .A1(b[11]), .A2(a[10]), .ZN(net215111) );
  XNOR2_X2 U8510 ( .A(net215211), .B(net215212), .ZN(net215209) );
  NAND2_X2 U8511 ( .A1(b[10]), .A2(a[11]), .ZN(n6081) );
  INV_X4 U8512 ( .A(n6081), .ZN(n6079) );
  NAND2_X2 U8513 ( .A1(b[9]), .A2(a[12]), .ZN(net215126) );
  NAND2_X2 U8514 ( .A1(b[8]), .A2(a[13]), .ZN(n6076) );
  INV_X4 U8515 ( .A(n6076), .ZN(n6073) );
  INV_X4 U8516 ( .A(net215206), .ZN(net215204) );
  NOR2_X4 U8517 ( .A1(net215204), .A2(n6022), .ZN(n6025) );
  INV_X4 U8518 ( .A(n6155), .ZN(n6027) );
  NAND3_X2 U8519 ( .A1(n5817), .A2(net215199), .A3(n6026), .ZN(n6153) );
  NAND2_X2 U8520 ( .A1(b[7]), .A2(a[14]), .ZN(n6068) );
  NAND2_X2 U8521 ( .A1(n6158), .A2(n6157), .ZN(n6066) );
  INV_X4 U8522 ( .A(n6030), .ZN(n6032) );
  NAND2_X2 U8523 ( .A1(n6163), .A2(n6162), .ZN(n6060) );
  NAND2_X2 U8524 ( .A1(net218536), .A2(a[18]), .ZN(n6042) );
  INV_X4 U8525 ( .A(net215175), .ZN(net215176) );
  NAND3_X4 U8526 ( .A1(net215176), .A2(a[19]), .A3(net218546), .ZN(n6173) );
  NAND2_X2 U8527 ( .A1(net218548), .A2(a[19]), .ZN(n6037) );
  NAND2_X2 U8528 ( .A1(n6037), .A2(net215175), .ZN(n6038) );
  NAND2_X2 U8529 ( .A1(n6173), .A2(n6038), .ZN(n6174) );
  XNOR2_X2 U8530 ( .A(n6172), .B(n6174), .ZN(n6039) );
  INV_X4 U8531 ( .A(n6039), .ZN(n6041) );
  INV_X4 U8532 ( .A(n6335), .ZN(n6040) );
  AOI21_X4 U8533 ( .B1(n6042), .B2(n6041), .A(n6040), .ZN(n6171) );
  INV_X4 U8534 ( .A(n6043), .ZN(n6046) );
  OAI21_X4 U8535 ( .B1(n6046), .B2(n6045), .A(n6044), .ZN(n6170) );
  INV_X4 U8536 ( .A(n6170), .ZN(n6047) );
  XNOR2_X2 U8537 ( .A(n6171), .B(n6047), .ZN(n6048) );
  INV_X4 U8538 ( .A(n6049), .ZN(n6052) );
  OAI21_X4 U8539 ( .B1(n6052), .B2(n6051), .A(n6050), .ZN(n6053) );
  INV_X4 U8540 ( .A(n6053), .ZN(n6169) );
  XNOR2_X2 U8541 ( .A(n6054), .B(n6169), .ZN(n6057) );
  INV_X4 U8542 ( .A(n6057), .ZN(n6055) );
  NAND2_X2 U8543 ( .A1(b[5]), .A2(a[16]), .ZN(n6056) );
  NAND2_X2 U8544 ( .A1(n6055), .A2(n6056), .ZN(n6164) );
  INV_X4 U8545 ( .A(n6056), .ZN(n6058) );
  NAND2_X2 U8546 ( .A1(n6058), .A2(n6057), .ZN(n6325) );
  XNOR2_X2 U8547 ( .A(n6060), .B(n6059), .ZN(n6063) );
  NAND2_X2 U8548 ( .A1(b[6]), .A2(a[15]), .ZN(n6062) );
  INV_X4 U8549 ( .A(n6062), .ZN(n6064) );
  NAND2_X2 U8550 ( .A1(n6064), .A2(n6063), .ZN(n6320) );
  XNOR2_X2 U8551 ( .A(n6066), .B(n6065), .ZN(n6069) );
  INV_X4 U8552 ( .A(n6069), .ZN(n6067) );
  INV_X4 U8553 ( .A(n6068), .ZN(n6070) );
  NAND2_X2 U8554 ( .A1(n6070), .A2(n6069), .ZN(n6315) );
  XNOR2_X2 U8555 ( .A(n6072), .B(n6071), .ZN(n6074) );
  NAND2_X2 U8556 ( .A1(n3904), .A2(n6073), .ZN(n6308) );
  INV_X4 U8557 ( .A(n6074), .ZN(n6075) );
  INV_X4 U8558 ( .A(n6077), .ZN(n6078) );
  XNOR2_X2 U8559 ( .A(net215129), .B(n6078), .ZN(net215127) );
  XNOR2_X2 U8560 ( .A(net215122), .B(net215121), .ZN(n6080) );
  NOR2_X4 U8561 ( .A1(n6307), .A2(n6082), .ZN(n6083) );
  XNOR2_X2 U8562 ( .A(net215114), .B(n6083), .ZN(net215112) );
  NAND2_X2 U8563 ( .A1(net214731), .A2(net214732), .ZN(n6084) );
  INV_X4 U8564 ( .A(net214804), .ZN(net214728) );
  AOI21_X4 U8565 ( .B1(n6084), .B2(net224078), .A(net214728), .ZN(n6085) );
  NAND2_X2 U8566 ( .A1(a[3]), .A2(b[18]), .ZN(net215062) );
  NAND2_X2 U8567 ( .A1(b[19]), .A2(a[2]), .ZN(n6252) );
  XNOR2_X2 U8568 ( .A(net215059), .B(n6252), .ZN(n6086) );
  XNOR2_X2 U8569 ( .A(n6086), .B(net219931), .ZN(n6430) );
  INV_X4 U8570 ( .A(n6088), .ZN(n6090) );
  NAND2_X2 U8571 ( .A1(n6426), .A2(n6428), .ZN(n6091) );
  NAND2_X2 U8572 ( .A1(b[20]), .A2(a[1]), .ZN(n6093) );
  INV_X4 U8573 ( .A(n6093), .ZN(n6096) );
  INV_X4 U8574 ( .A(n6094), .ZN(n6095) );
  NAND2_X2 U8575 ( .A1(n6101), .A2(n7805), .ZN(n6452) );
  OAI22_X2 U8576 ( .A1(n5042), .A2(n6452), .B1(n6102), .B2(n6454), .ZN(n6103)
         );
  NOR3_X4 U8577 ( .A1(n6104), .A2(n6103), .A3(n6639), .ZN(n6130) );
  INV_X4 U8578 ( .A(a[21]), .ZN(net215014) );
  INV_X4 U8579 ( .A(n6105), .ZN(n6106) );
  AOI22_X2 U8580 ( .A1(n6107), .A2(n3335), .B1(a[20]), .B2(n6106), .ZN(n6142)
         );
  XNOR2_X2 U8581 ( .A(n4002), .B(b[21]), .ZN(n6143) );
  XNOR2_X2 U8582 ( .A(n6143), .B(net215014), .ZN(n6141) );
  XNOR2_X2 U8583 ( .A(n6142), .B(n6141), .ZN(n6111) );
  INV_X4 U8584 ( .A(n6108), .ZN(n6109) );
  NAND2_X2 U8585 ( .A1(net218639), .A2(n6109), .ZN(n6110) );
  OAI221_X2 U8586 ( .B1(net215014), .B2(net218610), .C1(n7389), .C2(n6111), 
        .A(n6110), .ZN(n6120) );
  NAND2_X2 U8587 ( .A1(n6468), .A2(n6112), .ZN(n6118) );
  NAND2_X2 U8588 ( .A1(n6851), .A2(n6849), .ZN(n6117) );
  NAND2_X2 U8589 ( .A1(n7040), .A2(n6113), .ZN(n6116) );
  NAND4_X2 U8590 ( .A1(net215022), .A2(net215023), .A3(net215024), .A4(n6114), 
        .ZN(n7222) );
  NAND2_X2 U8591 ( .A1(n7050), .A2(n7222), .ZN(n6115) );
  NAND4_X2 U8592 ( .A1(n6118), .A2(n6117), .A3(n6116), .A4(n6115), .ZN(n6119)
         );
  NOR2_X4 U8593 ( .A1(n6120), .A2(n6119), .ZN(n6129) );
  INV_X4 U8594 ( .A(n6121), .ZN(n6269) );
  OAI221_X2 U8595 ( .B1(net215014), .B2(net218600), .C1(n6269), .C2(n7888), 
        .A(net218610), .ZN(n6127) );
  INV_X4 U8596 ( .A(n6850), .ZN(n6122) );
  INV_X4 U8597 ( .A(n6123), .ZN(n6124) );
  AOI211_X4 U8598 ( .C1(b[21]), .C2(n6127), .A(n6126), .B(n6125), .ZN(n6128)
         );
  INV_X4 U8599 ( .A(n6131), .ZN(n6136) );
  NOR2_X4 U8600 ( .A1(n6132), .A2(n3368), .ZN(n6134) );
  MUX2_X2 U8601 ( .A(net214224), .B(net215001), .S(net218558), .Z(n6133) );
  NAND2_X2 U8602 ( .A1(n6134), .A2(n6133), .ZN(n7802) );
  INV_X4 U8603 ( .A(n7802), .ZN(n6981) );
  OAI22_X2 U8604 ( .A1(n6136), .A2(n6637), .B1(n6981), .B2(n6135), .ZN(n6140)
         );
  INV_X4 U8605 ( .A(n6137), .ZN(n6138) );
  INV_X4 U8606 ( .A(n7806), .ZN(n6985) );
  OAI22_X2 U8607 ( .A1(n6138), .A2(n7035), .B1(n6985), .B2(n7053), .ZN(n6139)
         );
  NOR2_X4 U8608 ( .A1(n6140), .A2(n6139), .ZN(n6286) );
  XNOR2_X2 U8609 ( .A(n4002), .B(b[22]), .ZN(n6459) );
  XNOR2_X2 U8610 ( .A(n6459), .B(net214758), .ZN(n6458) );
  OAI22_X2 U8611 ( .A1(n6143), .A2(net215014), .B1(n6142), .B2(n6141), .ZN(
        n6462) );
  XNOR2_X2 U8612 ( .A(n6458), .B(n6462), .ZN(n6147) );
  AOI211_X4 U8613 ( .C1(n6147), .C2(n3990), .A(n6146), .B(n6145), .ZN(n6285)
         );
  NAND2_X2 U8614 ( .A1(net218658), .A2(net214984), .ZN(n6271) );
  NAND2_X2 U8615 ( .A1(b[16]), .A2(a[6]), .ZN(n6247) );
  INV_X4 U8616 ( .A(n6247), .ZN(n6246) );
  NAND2_X2 U8617 ( .A1(b[15]), .A2(a[7]), .ZN(n6241) );
  INV_X4 U8618 ( .A(n6241), .ZN(n6240) );
  AOI21_X4 U8619 ( .B1(n3941), .B2(n6149), .A(net214978), .ZN(net214974) );
  OAI21_X4 U8620 ( .B1(net214963), .B2(net214964), .A(n6150), .ZN(n6305) );
  NAND2_X2 U8621 ( .A1(a[13]), .A2(b[9]), .ZN(n6215) );
  INV_X4 U8622 ( .A(n6215), .ZN(n6212) );
  NAND2_X2 U8623 ( .A1(n6309), .A2(n6308), .ZN(n6211) );
  NAND2_X2 U8624 ( .A1(b[8]), .A2(a[14]), .ZN(n6209) );
  INV_X4 U8625 ( .A(n6209), .ZN(n6206) );
  INV_X4 U8626 ( .A(n6153), .ZN(n6156) );
  OAI21_X4 U8627 ( .B1(n6156), .B2(n6155), .A(n6154), .ZN(n6316) );
  NAND2_X2 U8628 ( .A1(n6316), .A2(n3905), .ZN(n6205) );
  INV_X4 U8629 ( .A(n6157), .ZN(n6161) );
  INV_X4 U8630 ( .A(n6158), .ZN(n6160) );
  OAI21_X4 U8631 ( .B1(n6161), .B2(n6160), .A(n6159), .ZN(n6321) );
  NAND2_X2 U8632 ( .A1(n6321), .A2(n6320), .ZN(n6199) );
  INV_X4 U8633 ( .A(n6162), .ZN(n6166) );
  INV_X4 U8634 ( .A(n6163), .ZN(n6165) );
  OAI21_X4 U8635 ( .B1(n6166), .B2(n6165), .A(n6164), .ZN(n6326) );
  NAND2_X2 U8636 ( .A1(a[18]), .A2(b[4]), .ZN(n6186) );
  INV_X4 U8637 ( .A(n6186), .ZN(n6183) );
  NAND2_X2 U8638 ( .A1(net218536), .A2(a[19]), .ZN(n6179) );
  OAI21_X4 U8639 ( .B1(n6175), .B2(n6174), .A(n6173), .ZN(n6341) );
  NAND3_X2 U8640 ( .A1(a[20]), .A2(net214922), .A3(net218548), .ZN(n6541) );
  NAND2_X2 U8641 ( .A1(net218548), .A2(a[20]), .ZN(n6176) );
  INV_X4 U8642 ( .A(net214922), .ZN(net214921) );
  NAND2_X2 U8643 ( .A1(n6176), .A2(net214921), .ZN(n6340) );
  NAND2_X2 U8644 ( .A1(n6541), .A2(n6340), .ZN(n6177) );
  XNOR2_X2 U8645 ( .A(n6341), .B(n6177), .ZN(n6180) );
  INV_X4 U8646 ( .A(n6180), .ZN(n6178) );
  NAND2_X2 U8647 ( .A1(n6179), .A2(n6178), .ZN(n6181) );
  NAND3_X2 U8648 ( .A1(a[19]), .A2(n6180), .A3(net218536), .ZN(n6337) );
  NAND2_X2 U8649 ( .A1(n6181), .A2(n6337), .ZN(n6338) );
  XNOR2_X2 U8650 ( .A(n6182), .B(n6338), .ZN(n6184) );
  NAND2_X2 U8651 ( .A1(n6183), .A2(n6184), .ZN(n6332) );
  INV_X4 U8652 ( .A(n6184), .ZN(n6185) );
  NAND2_X2 U8653 ( .A1(n6186), .A2(n6185), .ZN(n6330) );
  NAND2_X2 U8654 ( .A1(n6332), .A2(n6330), .ZN(n6187) );
  XNOR2_X2 U8655 ( .A(n6331), .B(n6187), .ZN(n6190) );
  INV_X4 U8656 ( .A(n6190), .ZN(n6188) );
  NAND2_X2 U8657 ( .A1(a[17]), .A2(b[5]), .ZN(n6189) );
  NAND2_X2 U8658 ( .A1(n6188), .A2(n6189), .ZN(n6327) );
  INV_X4 U8659 ( .A(n6189), .ZN(n6191) );
  NAND2_X2 U8660 ( .A1(n6191), .A2(n6190), .ZN(n6527) );
  NAND2_X2 U8661 ( .A1(n6327), .A2(n6527), .ZN(n6192) );
  XNOR2_X2 U8662 ( .A(n6193), .B(n6192), .ZN(n6196) );
  NAND2_X2 U8663 ( .A1(a[16]), .A2(b[6]), .ZN(n6195) );
  INV_X4 U8664 ( .A(n6195), .ZN(n6197) );
  XNOR2_X2 U8665 ( .A(n6199), .B(n6198), .ZN(n6202) );
  INV_X4 U8666 ( .A(n6202), .ZN(n6200) );
  NAND2_X2 U8667 ( .A1(b[7]), .A2(a[15]), .ZN(n6201) );
  NAND2_X2 U8668 ( .A1(n6200), .A2(n6201), .ZN(n6317) );
  INV_X4 U8669 ( .A(n6201), .ZN(n6203) );
  NAND2_X2 U8670 ( .A1(n6203), .A2(n6202), .ZN(n6514) );
  NAND2_X2 U8671 ( .A1(n6317), .A2(n6514), .ZN(n6204) );
  XNOR2_X2 U8672 ( .A(n6205), .B(n6204), .ZN(n6207) );
  NAND2_X2 U8673 ( .A1(n6206), .A2(n6207), .ZN(n6313) );
  INV_X4 U8674 ( .A(n6207), .ZN(n6208) );
  XNOR2_X2 U8675 ( .A(n6211), .B(n6210), .ZN(n6213) );
  NAND2_X2 U8676 ( .A1(n6212), .A2(n6213), .ZN(net214429) );
  INV_X4 U8677 ( .A(net214429), .ZN(net214620) );
  NOR2_X4 U8678 ( .A1(net214620), .A2(net214427), .ZN(n6216) );
  XNOR2_X2 U8679 ( .A(n6216), .B(net214428), .ZN(n6219) );
  INV_X4 U8680 ( .A(n6219), .ZN(n6217) );
  NAND2_X2 U8681 ( .A1(a[12]), .A2(b[10]), .ZN(n6218) );
  INV_X4 U8682 ( .A(n6218), .ZN(n6220) );
  INV_X4 U8683 ( .A(n6229), .ZN(n6225) );
  NAND2_X2 U8684 ( .A1(b[12]), .A2(a[10]), .ZN(n6227) );
  OAI21_X4 U8685 ( .B1(n6226), .B2(n6225), .A(n6227), .ZN(n6303) );
  INV_X4 U8686 ( .A(n6227), .ZN(n6228) );
  XNOR2_X2 U8687 ( .A(n6230), .B(n6302), .ZN(n6232) );
  NAND2_X2 U8688 ( .A1(b[13]), .A2(a[9]), .ZN(n6231) );
  INV_X4 U8689 ( .A(n6231), .ZN(n6233) );
  NAND2_X2 U8690 ( .A1(b[14]), .A2(a[8]), .ZN(n6235) );
  NAND2_X2 U8691 ( .A1(n6235), .A2(n6236), .ZN(n6301) );
  INV_X4 U8692 ( .A(n6235), .ZN(n6238) );
  NAND2_X2 U8693 ( .A1(n3790), .A2(n6240), .ZN(n6410) );
  INV_X4 U8694 ( .A(n3940), .ZN(n6242) );
  XNOR2_X2 U8695 ( .A(net214792), .B(net214793), .ZN(n6250) );
  NAND2_X2 U8696 ( .A1(a[3]), .A2(b[19]), .ZN(n6249) );
  INV_X4 U8697 ( .A(n6249), .ZN(n6251) );
  NAND2_X2 U8698 ( .A1(n6251), .A2(n6250), .ZN(n6432) );
  NAND2_X2 U8699 ( .A1(n6425), .A2(n6432), .ZN(n6257) );
  INV_X4 U8700 ( .A(n6252), .ZN(n6254) );
  XNOR2_X2 U8701 ( .A(net214784), .B(net214785), .ZN(n6253) );
  NAND2_X2 U8702 ( .A1(n6255), .A2(n6427), .ZN(n6256) );
  XNOR2_X2 U8703 ( .A(n6257), .B(n6256), .ZN(n6260) );
  INV_X4 U8704 ( .A(n6260), .ZN(n6258) );
  NAND2_X2 U8705 ( .A1(b[20]), .A2(a[2]), .ZN(n6259) );
  INV_X4 U8706 ( .A(n6259), .ZN(n6261) );
  NAND2_X2 U8707 ( .A1(n6261), .A2(n6260), .ZN(n6297) );
  INV_X4 U8708 ( .A(n6295), .ZN(n6262) );
  XNOR2_X2 U8709 ( .A(n6263), .B(n6264), .ZN(n6267) );
  INV_X4 U8710 ( .A(n6267), .ZN(n6265) );
  NAND2_X2 U8711 ( .A1(b[21]), .A2(a[1]), .ZN(n6266) );
  NAND2_X2 U8712 ( .A1(n6265), .A2(n6266), .ZN(n6287) );
  INV_X4 U8713 ( .A(n6266), .ZN(n6268) );
  NAND2_X2 U8714 ( .A1(n6268), .A2(n6267), .ZN(n6288) );
  NAND3_X4 U8715 ( .A1(a[0]), .A2(b[21]), .A3(n6269), .ZN(n6289) );
  XNOR2_X2 U8716 ( .A(n6270), .B(n6289), .ZN(n6276) );
  OAI22_X2 U8717 ( .A1(n4766), .A2(n6452), .B1(n6273), .B2(n6454), .ZN(n6274)
         );
  NOR3_X4 U8718 ( .A1(n6275), .A2(n6274), .A3(n6639), .ZN(n6284) );
  INV_X4 U8719 ( .A(n6276), .ZN(n6447) );
  OAI221_X2 U8720 ( .B1(net214758), .B2(net218600), .C1(n6447), .C2(net218655), 
        .A(net218610), .ZN(n6282) );
  INV_X4 U8721 ( .A(n6278), .ZN(n6279) );
  AOI211_X4 U8722 ( .C1(b[22]), .C2(n6282), .A(n6281), .B(n6280), .ZN(n6283)
         );
  NAND4_X2 U8723 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(
        result[22]) );
  NAND2_X2 U8724 ( .A1(net218658), .A2(net214747), .ZN(n6450) );
  OAI21_X4 U8725 ( .B1(n6290), .B2(n6289), .A(n6288), .ZN(n6441) );
  INV_X4 U8726 ( .A(n6291), .ZN(n6299) );
  AOI21_X4 U8727 ( .B1(n6296), .B2(n6295), .A(n6294), .ZN(n6298) );
  OAI21_X4 U8728 ( .B1(n6299), .B2(n6298), .A(n6297), .ZN(n6609) );
  XNOR2_X2 U8729 ( .A(n6676), .B(n3376), .ZN(n6440) );
  NAND2_X2 U8730 ( .A1(b[17]), .A2(a[6]), .ZN(n6421) );
  INV_X4 U8731 ( .A(n6421), .ZN(n6419) );
  NAND2_X2 U8732 ( .A1(b[16]), .A2(a[7]), .ZN(n6415) );
  INV_X4 U8733 ( .A(n6415), .ZN(n6413) );
  NAND2_X2 U8734 ( .A1(n6494), .A2(n6493), .ZN(n6404) );
  NAND2_X2 U8735 ( .A1(b[14]), .A2(a[9]), .ZN(n6401) );
  INV_X4 U8736 ( .A(n6401), .ZN(n6399) );
  INV_X4 U8737 ( .A(n6302), .ZN(n6304) );
  NAND2_X2 U8738 ( .A1(b[12]), .A2(a[11]), .ZN(n6389) );
  INV_X4 U8739 ( .A(n6389), .ZN(n6387) );
  OAI21_X4 U8740 ( .B1(n6306), .B2(n6307), .A(net214705), .ZN(net214433) );
  NAND2_X2 U8741 ( .A1(a[13]), .A2(b[10]), .ZN(net214612) );
  NAND2_X2 U8742 ( .A1(a[14]), .A2(b[9]), .ZN(n6375) );
  INV_X4 U8743 ( .A(n6308), .ZN(n6312) );
  INV_X4 U8744 ( .A(n6309), .ZN(n6311) );
  OAI21_X4 U8745 ( .B1(n6312), .B2(n6311), .A(n6310), .ZN(n6314) );
  INV_X4 U8746 ( .A(n6316), .ZN(n6318) );
  OAI21_X4 U8747 ( .B1(n6319), .B2(n6318), .A(n6317), .ZN(n6515) );
  INV_X4 U8748 ( .A(n6321), .ZN(n6323) );
  OAI21_X4 U8749 ( .B1(n6324), .B2(n6323), .A(n6322), .ZN(n6520) );
  INV_X4 U8750 ( .A(n6326), .ZN(n6328) );
  OAI21_X4 U8751 ( .B1(n6329), .B2(n6328), .A(n6327), .ZN(n6526) );
  NAND2_X2 U8752 ( .A1(n6526), .A2(n6527), .ZN(n6356) );
  NAND2_X2 U8753 ( .A1(a[18]), .A2(b[5]), .ZN(n6354) );
  INV_X4 U8754 ( .A(n6354), .ZN(n6351) );
  NAND2_X2 U8755 ( .A1(n6331), .A2(n6330), .ZN(n6333) );
  INV_X4 U8756 ( .A(n6336), .ZN(n6339) );
  OAI21_X4 U8757 ( .B1(n6339), .B2(n6338), .A(n6337), .ZN(n6536) );
  NAND2_X2 U8758 ( .A1(net218536), .A2(a[20]), .ZN(n6346) );
  NAND2_X2 U8759 ( .A1(n6341), .A2(n6340), .ZN(n6542) );
  INV_X4 U8760 ( .A(net214660), .ZN(net214661) );
  NAND3_X4 U8761 ( .A1(net214661), .A2(a[21]), .A3(net218546), .ZN(n6543) );
  NAND2_X2 U8762 ( .A1(net218548), .A2(a[21]), .ZN(n6342) );
  NAND2_X2 U8763 ( .A1(n6342), .A2(net214660), .ZN(n6545) );
  NAND2_X2 U8764 ( .A1(n6543), .A2(n6545), .ZN(n6343) );
  XNOR2_X2 U8765 ( .A(n6344), .B(n6343), .ZN(n6347) );
  INV_X4 U8766 ( .A(n6347), .ZN(n6345) );
  NAND2_X2 U8767 ( .A1(n6346), .A2(n6345), .ZN(n6348) );
  NAND3_X2 U8768 ( .A1(a[20]), .A2(n6347), .A3(net218534), .ZN(n6537) );
  XNOR2_X2 U8769 ( .A(n6536), .B(n6538), .ZN(n6349) );
  NAND3_X2 U8770 ( .A1(a[19]), .A2(n6349), .A3(b[4]), .ZN(n6534) );
  XNOR2_X2 U8771 ( .A(n6533), .B(n6350), .ZN(n6352) );
  NAND2_X2 U8772 ( .A1(n6351), .A2(n6352), .ZN(n6528) );
  INV_X4 U8773 ( .A(n6352), .ZN(n6353) );
  NAND2_X2 U8774 ( .A1(n6354), .A2(n6353), .ZN(n6531) );
  NAND2_X2 U8775 ( .A1(n6528), .A2(n6531), .ZN(n6355) );
  XNOR2_X2 U8776 ( .A(n6356), .B(n6355), .ZN(n6359) );
  INV_X4 U8777 ( .A(n6359), .ZN(n6357) );
  NAND2_X2 U8778 ( .A1(a[17]), .A2(b[6]), .ZN(n6358) );
  NAND2_X2 U8779 ( .A1(n6357), .A2(n6358), .ZN(n6521) );
  INV_X4 U8780 ( .A(n6358), .ZN(n6360) );
  NAND2_X2 U8781 ( .A1(n6360), .A2(n6359), .ZN(n6524) );
  NAND2_X2 U8782 ( .A1(n6521), .A2(n6524), .ZN(n6361) );
  XNOR2_X2 U8783 ( .A(n6362), .B(n6361), .ZN(n6365) );
  INV_X4 U8784 ( .A(n6365), .ZN(n6363) );
  NAND2_X2 U8785 ( .A1(b[7]), .A2(a[16]), .ZN(n6364) );
  NAND2_X2 U8786 ( .A1(n6363), .A2(n6364), .ZN(n6516) );
  INV_X4 U8787 ( .A(n6364), .ZN(n6366) );
  XNOR2_X2 U8788 ( .A(n6368), .B(n6367), .ZN(n6371) );
  INV_X4 U8789 ( .A(n6371), .ZN(n6369) );
  NAND2_X2 U8790 ( .A1(b[8]), .A2(a[15]), .ZN(n6370) );
  INV_X4 U8791 ( .A(n6370), .ZN(n6372) );
  XNOR2_X2 U8792 ( .A(n6513), .B(n6373), .ZN(n6376) );
  INV_X4 U8793 ( .A(n6376), .ZN(n6374) );
  NAND2_X2 U8794 ( .A1(n6375), .A2(n6374), .ZN(n6510) );
  INV_X4 U8795 ( .A(n6375), .ZN(n6377) );
  NAND2_X2 U8796 ( .A1(a[12]), .A2(b[11]), .ZN(n6380) );
  INV_X4 U8797 ( .A(n6380), .ZN(n6381) );
  NAND2_X2 U8798 ( .A1(n3590), .A2(n6384), .ZN(n6507) );
  XNOR2_X2 U8799 ( .A(n6386), .B(n6385), .ZN(n6388) );
  NAND2_X2 U8800 ( .A1(n6387), .A2(n6388), .ZN(n6504) );
  INV_X4 U8801 ( .A(n6388), .ZN(n6390) );
  XNOR2_X2 U8802 ( .A(n6391), .B(n6392), .ZN(n6395) );
  INV_X4 U8803 ( .A(n6395), .ZN(n6393) );
  NAND2_X2 U8804 ( .A1(b[13]), .A2(a[10]), .ZN(n6394) );
  INV_X4 U8805 ( .A(n6394), .ZN(n6396) );
  OAI21_X4 U8806 ( .B1(net214583), .B2(net214584), .A(n6397), .ZN(n6708) );
  XNOR2_X2 U8807 ( .A(n6398), .B(n6708), .ZN(n6400) );
  XNOR2_X2 U8808 ( .A(n6404), .B(n6403), .ZN(n6407) );
  NAND2_X2 U8809 ( .A1(b[15]), .A2(a[8]), .ZN(n6406) );
  INV_X4 U8810 ( .A(n6406), .ZN(n6408) );
  XNOR2_X2 U8811 ( .A(n6412), .B(n6693), .ZN(n6414) );
  XNOR2_X2 U8812 ( .A(n6417), .B(n6418), .ZN(n6420) );
  INV_X4 U8813 ( .A(n3426), .ZN(n6422) );
  NAND2_X2 U8814 ( .A1(b[19]), .A2(net219055), .ZN(n6423) );
  INV_X4 U8815 ( .A(n6423), .ZN(n6424) );
  NAND2_X2 U8816 ( .A1(n6424), .A2(net214536), .ZN(n6685) );
  INV_X4 U8817 ( .A(n6425), .ZN(n6434) );
  NAND3_X2 U8818 ( .A1(n6426), .A2(n6427), .A3(n6428), .ZN(n6429) );
  OAI21_X4 U8819 ( .B1(n6433), .B2(n6434), .A(n6432), .ZN(n6680) );
  XNOR2_X2 U8820 ( .A(n6680), .B(n6435), .ZN(n6438) );
  INV_X4 U8821 ( .A(n6438), .ZN(n6436) );
  NAND2_X2 U8822 ( .A1(a[3]), .A2(b[20]), .ZN(n6437) );
  INV_X4 U8823 ( .A(n6437), .ZN(n6439) );
  NAND2_X2 U8824 ( .A1(n6439), .A2(n6438), .ZN(n6675) );
  NAND2_X2 U8825 ( .A1(n6674), .A2(n6675), .ZN(n6610) );
  XNOR2_X2 U8826 ( .A(n6440), .B(n6610), .ZN(n6442) );
  INV_X4 U8827 ( .A(n6442), .ZN(n6668) );
  NAND2_X2 U8828 ( .A1(n6669), .A2(n6668), .ZN(n6443) );
  NAND2_X2 U8829 ( .A1(n6442), .A2(n6441), .ZN(n6612) );
  NAND2_X2 U8830 ( .A1(n6443), .A2(n6612), .ZN(n6446) );
  INV_X4 U8831 ( .A(n6445), .ZN(n6486) );
  INV_X4 U8832 ( .A(n6446), .ZN(n6485) );
  INV_X4 U8833 ( .A(n6664), .ZN(n6444) );
  NAND3_X4 U8834 ( .A1(b[22]), .A2(a[0]), .A3(n6447), .ZN(n6483) );
  XNOR2_X2 U8835 ( .A(n6448), .B(n6483), .ZN(n6625) );
  INV_X4 U8836 ( .A(n6451), .ZN(n6455) );
  OAI22_X2 U8837 ( .A1(n6455), .A2(n6454), .B1(n6453), .B2(n6452), .ZN(n6456)
         );
  NOR3_X4 U8838 ( .A1(n6457), .A2(n6456), .A3(n6639), .ZN(n6482) );
  INV_X4 U8839 ( .A(a[23]), .ZN(net214479) );
  INV_X4 U8840 ( .A(n6458), .ZN(n6461) );
  INV_X4 U8841 ( .A(n6459), .ZN(n6460) );
  AOI22_X2 U8842 ( .A1(n6462), .A2(n6461), .B1(a[22]), .B2(n6460), .ZN(n6643)
         );
  XNOR2_X2 U8843 ( .A(n4002), .B(b[23]), .ZN(n6644) );
  XNOR2_X2 U8844 ( .A(n6644), .B(net214479), .ZN(n6642) );
  XNOR2_X2 U8845 ( .A(n6643), .B(n6642), .ZN(n6466) );
  INV_X4 U8846 ( .A(n6463), .ZN(n6464) );
  NAND2_X2 U8847 ( .A1(net218639), .A2(n6464), .ZN(n6465) );
  OAI221_X2 U8848 ( .B1(net214479), .B2(net218610), .C1(n7389), .C2(n6466), 
        .A(n6465), .ZN(n6476) );
  NAND2_X2 U8849 ( .A1(n6468), .A2(n6467), .ZN(n6474) );
  NAND2_X2 U8850 ( .A1(n6851), .A2(net212010), .ZN(n6473) );
  NAND2_X2 U8851 ( .A1(n7040), .A2(n6469), .ZN(n6472) );
  NAND4_X2 U8852 ( .A1(net214486), .A2(net214487), .A3(n6470), .A4(net214489), 
        .ZN(n7046) );
  NAND2_X2 U8853 ( .A1(n7050), .A2(n7046), .ZN(n6471) );
  NAND4_X2 U8854 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6475)
         );
  NOR2_X4 U8855 ( .A1(n6476), .A2(n6475), .ZN(n6481) );
  INV_X4 U8856 ( .A(net213359), .ZN(net214478) );
  INV_X4 U8857 ( .A(net214477), .ZN(net214476) );
  INV_X4 U8858 ( .A(n6483), .ZN(n6484) );
  OAI21_X4 U8859 ( .B1(n6486), .B2(n6485), .A(n6484), .ZN(n6665) );
  INV_X4 U8860 ( .A(n6681), .ZN(n6488) );
  OAI21_X4 U8861 ( .B1(n6488), .B2(n6487), .A(n3967), .ZN(n6600) );
  NAND2_X2 U8862 ( .A1(b[18]), .A2(a[6]), .ZN(net214293) );
  INV_X4 U8863 ( .A(n6694), .ZN(n6492) );
  INV_X4 U8864 ( .A(n6693), .ZN(n6491) );
  OAI21_X4 U8865 ( .B1(n6491), .B2(n6492), .A(n6697), .ZN(n6585) );
  NAND2_X2 U8866 ( .A1(n6494), .A2(n6493), .ZN(n6496) );
  INV_X4 U8867 ( .A(n6708), .ZN(n6497) );
  INV_X4 U8868 ( .A(n6499), .ZN(n6503) );
  INV_X4 U8869 ( .A(n6500), .ZN(n6502) );
  OAI21_X4 U8870 ( .B1(n6503), .B2(n6502), .A(n6501), .ZN(n6505) );
  INV_X4 U8871 ( .A(n6713), .ZN(n6508) );
  OAI21_X4 U8872 ( .B1(n6509), .B2(n6508), .A(n6710), .ZN(net213557) );
  NAND2_X2 U8873 ( .A1(a[13]), .A2(b[11]), .ZN(net214331) );
  INV_X4 U8874 ( .A(net214331), .ZN(net214334) );
  NAND2_X2 U8875 ( .A1(n6511), .A2(n6510), .ZN(n6716) );
  NAND2_X2 U8876 ( .A1(n6716), .A2(n6715), .ZN(n6573) );
  NAND2_X2 U8877 ( .A1(n6513), .A2(n6512), .ZN(n6721) );
  INV_X4 U8878 ( .A(n6515), .ZN(n6517) );
  OAI21_X4 U8879 ( .B1(n6518), .B2(n6517), .A(n6516), .ZN(n6727) );
  NAND2_X2 U8880 ( .A1(n6727), .A2(n6726), .ZN(n6563) );
  INV_X4 U8881 ( .A(n6520), .ZN(n6522) );
  NAND2_X2 U8882 ( .A1(n6525), .A2(n6524), .ZN(n6734) );
  NAND2_X2 U8883 ( .A1(a[18]), .A2(b[6]), .ZN(n6556) );
  INV_X4 U8884 ( .A(n6556), .ZN(n6554) );
  NAND2_X2 U8885 ( .A1(n6527), .A2(n6526), .ZN(n6530) );
  INV_X4 U8886 ( .A(n6528), .ZN(n6529) );
  AOI21_X4 U8887 ( .B1(n6531), .B2(n6530), .A(n6529), .ZN(n6740) );
  NAND2_X2 U8888 ( .A1(a[19]), .A2(b[5]), .ZN(n6552) );
  INV_X4 U8889 ( .A(n6552), .ZN(n6549) );
  INV_X4 U8890 ( .A(n6533), .ZN(n6535) );
  OAI21_X4 U8891 ( .B1(n3758), .B2(n6535), .A(n6534), .ZN(n6742) );
  INV_X4 U8892 ( .A(n6536), .ZN(n6539) );
  OAI21_X4 U8893 ( .B1(n6539), .B2(n6538), .A(n6537), .ZN(net214084) );
  NAND2_X2 U8894 ( .A1(a[22]), .A2(net218550), .ZN(n6540) );
  NAND2_X2 U8895 ( .A1(n6540), .A2(net214387), .ZN(net214384) );
  INV_X4 U8896 ( .A(n6543), .ZN(n6544) );
  AOI21_X4 U8897 ( .B1(n6344), .B2(n6545), .A(n6544), .ZN(net214101) );
  NAND3_X2 U8898 ( .A1(a[21]), .A2(net214376), .A3(net218534), .ZN(net214083)
         );
  NAND2_X2 U8899 ( .A1(net218536), .A2(a[21]), .ZN(n6546) );
  NAND2_X2 U8900 ( .A1(n6546), .A2(net220496), .ZN(net214085) );
  NAND3_X2 U8901 ( .A1(a[20]), .A2(net214372), .A3(b[4]), .ZN(n6743) );
  NAND2_X2 U8902 ( .A1(a[20]), .A2(b[4]), .ZN(n6547) );
  INV_X4 U8903 ( .A(net214372), .ZN(net214371) );
  NAND2_X2 U8904 ( .A1(n6547), .A2(net214371), .ZN(n6548) );
  XNOR2_X2 U8905 ( .A(n6742), .B(n6744), .ZN(n6550) );
  NAND2_X2 U8906 ( .A1(n6549), .A2(n6550), .ZN(n6739) );
  INV_X4 U8907 ( .A(n6550), .ZN(n6551) );
  NAND2_X2 U8908 ( .A1(n6739), .A2(n6738), .ZN(n6553) );
  NAND2_X2 U8909 ( .A1(n6554), .A2(n6555), .ZN(n6735) );
  NAND2_X2 U8910 ( .A1(n6556), .A2(n3761), .ZN(n6733) );
  NAND2_X2 U8911 ( .A1(n6735), .A2(n6733), .ZN(n6557) );
  XNOR2_X2 U8912 ( .A(n6734), .B(n6557), .ZN(n6560) );
  INV_X4 U8913 ( .A(n6560), .ZN(n6558) );
  NAND2_X2 U8914 ( .A1(b[7]), .A2(a[17]), .ZN(n6559) );
  INV_X4 U8915 ( .A(n6559), .ZN(n6561) );
  NAND2_X2 U8916 ( .A1(n6561), .A2(n6560), .ZN(n6731) );
  XNOR2_X2 U8917 ( .A(n6563), .B(n6562), .ZN(n6724) );
  INV_X4 U8918 ( .A(n6724), .ZN(n6564) );
  NAND2_X2 U8919 ( .A1(b[8]), .A2(a[16]), .ZN(n6565) );
  INV_X4 U8920 ( .A(n6565), .ZN(n6725) );
  NAND2_X2 U8921 ( .A1(n6722), .A2(n6566), .ZN(n6567) );
  XNOR2_X2 U8922 ( .A(n6723), .B(n6567), .ZN(n6570) );
  INV_X4 U8923 ( .A(n6570), .ZN(n6568) );
  NAND2_X2 U8924 ( .A1(a[15]), .A2(b[9]), .ZN(n6569) );
  NAND2_X2 U8925 ( .A1(n6568), .A2(n6569), .ZN(n6717) );
  INV_X4 U8926 ( .A(n6569), .ZN(n6571) );
  NAND2_X2 U8927 ( .A1(n6571), .A2(n6570), .ZN(n6901) );
  XNOR2_X2 U8928 ( .A(n6573), .B(n6572), .ZN(net214338) );
  NAND2_X2 U8929 ( .A1(a[14]), .A2(b[10]), .ZN(net214339) );
  XNOR2_X2 U8930 ( .A(net214329), .B(net214330), .ZN(n6787) );
  INV_X4 U8931 ( .A(net214323), .ZN(net214326) );
  NAND2_X2 U8932 ( .A1(b[13]), .A2(a[11]), .ZN(net214325) );
  INV_X4 U8933 ( .A(net214325), .ZN(net214324) );
  XNOR2_X2 U8934 ( .A(n6577), .B(n6576), .ZN(n6580) );
  NAND2_X2 U8935 ( .A1(b[14]), .A2(a[10]), .ZN(n6579) );
  INV_X4 U8936 ( .A(n6579), .ZN(n6581) );
  NAND2_X2 U8937 ( .A1(n6581), .A2(n6580), .ZN(n6701) );
  XNOR2_X2 U8938 ( .A(n6704), .B(n6582), .ZN(n6583) );
  XNOR2_X2 U8939 ( .A(n6584), .B(n6585), .ZN(n6588) );
  NAND2_X2 U8940 ( .A1(b[16]), .A2(a[8]), .ZN(n6587) );
  INV_X4 U8941 ( .A(n6587), .ZN(n6589) );
  NAND2_X2 U8942 ( .A1(n6589), .A2(n3792), .ZN(n6691) );
  XNOR2_X2 U8943 ( .A(n6690), .B(n6590), .ZN(n6593) );
  INV_X4 U8944 ( .A(n3951), .ZN(n6591) );
  NAND2_X2 U8945 ( .A1(b[17]), .A2(a[7]), .ZN(n6592) );
  INV_X4 U8946 ( .A(n6592), .ZN(n6594) );
  XNOR2_X2 U8947 ( .A(net214288), .B(net214289), .ZN(n6597) );
  INV_X4 U8948 ( .A(n6597), .ZN(n6595) );
  NAND2_X2 U8949 ( .A1(b[19]), .A2(a[5]), .ZN(n6596) );
  INV_X4 U8950 ( .A(n6596), .ZN(n6598) );
  NAND2_X2 U8951 ( .A1(n6598), .A2(n6597), .ZN(n6878) );
  XNOR2_X2 U8952 ( .A(n6600), .B(n6599), .ZN(n6603) );
  NAND2_X2 U8953 ( .A1(b[20]), .A2(net219055), .ZN(n6602) );
  INV_X4 U8954 ( .A(n6602), .ZN(n6604) );
  NAND2_X2 U8955 ( .A1(n6604), .A2(n6603), .ZN(n6939) );
  XNOR2_X2 U8956 ( .A(n6606), .B(n6605), .ZN(n6670) );
  INV_X4 U8957 ( .A(n3911), .ZN(n6607) );
  NAND2_X2 U8958 ( .A1(a[3]), .A2(b[21]), .ZN(n6608) );
  INV_X4 U8959 ( .A(n6608), .ZN(n6671) );
  XNOR2_X2 U8960 ( .A(n6614), .B(n6613), .ZN(n6617) );
  INV_X4 U8961 ( .A(n3765), .ZN(n6615) );
  NAND2_X2 U8962 ( .A1(b[22]), .A2(a[2]), .ZN(n6616) );
  INV_X4 U8963 ( .A(n6616), .ZN(n6618) );
  NAND2_X2 U8964 ( .A1(n6666), .A2(n6955), .ZN(n6619) );
  XNOR2_X2 U8965 ( .A(n6620), .B(n6619), .ZN(n6623) );
  INV_X4 U8966 ( .A(n6623), .ZN(n6621) );
  NAND2_X2 U8967 ( .A1(b[23]), .A2(a[1]), .ZN(n6622) );
  INV_X4 U8968 ( .A(n6622), .ZN(n6624) );
  NAND2_X2 U8969 ( .A1(n6662), .A2(n6833), .ZN(n6626) );
  INV_X4 U8970 ( .A(n6627), .ZN(n6840) );
  AOI21_X2 U8971 ( .B1(b[24]), .B2(n6629), .A(n6628), .ZN(n6660) );
  NAND2_X2 U8972 ( .A1(n7033), .A2(n6630), .ZN(n6659) );
  NAND2_X2 U8973 ( .A1(net218658), .A2(net214247), .ZN(n6631) );
  NAND2_X2 U8974 ( .A1(n6631), .A2(net212094), .ZN(n6641) );
  XNOR2_X2 U8975 ( .A(n4002), .B(b[24]), .ZN(n6852) );
  OAI22_X2 U8976 ( .A1(n6644), .A2(net214479), .B1(n6643), .B2(n6642), .ZN(
        n6854) );
  XNOR2_X2 U8977 ( .A(n3336), .B(n6854), .ZN(n6649) );
  MUX2_X2 U8978 ( .A(net213634), .B(net214224), .S(net218558), .Z(n6646) );
  NAND2_X2 U8979 ( .A1(n6647), .A2(n6646), .ZN(n7073) );
  NAND2_X2 U8980 ( .A1(n7050), .A2(n7073), .ZN(n6648) );
  OAI221_X2 U8981 ( .B1(n3364), .B2(n7053), .C1(n7389), .C2(n6649), .A(n6648), 
        .ZN(n6656) );
  NAND2_X2 U8982 ( .A1(net218639), .A2(n6650), .ZN(n6651) );
  NOR3_X2 U8983 ( .A1(n6656), .A2(n6655), .A3(n6654), .ZN(n6657) );
  NAND4_X2 U8984 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(
        result[24]) );
  INV_X4 U8985 ( .A(n6661), .ZN(n6663) );
  NAND2_X2 U8986 ( .A1(b[23]), .A2(a[2]), .ZN(n6954) );
  XNOR2_X2 U8987 ( .A(n6954), .B(net213680), .ZN(n6830) );
  NAND2_X2 U8988 ( .A1(b[22]), .A2(a[3]), .ZN(n6828) );
  INV_X4 U8989 ( .A(n6828), .ZN(n6825) );
  OAI21_X4 U8990 ( .B1(n6669), .B2(n6668), .A(n6667), .ZN(n6872) );
  INV_X4 U8991 ( .A(n6876), .ZN(n6672) );
  OAI21_X4 U8992 ( .B1(n6673), .B2(n6672), .A(n6873), .ZN(n6824) );
  NAND2_X2 U8993 ( .A1(b[21]), .A2(net219055), .ZN(n6821) );
  INV_X4 U8994 ( .A(n6821), .ZN(n6819) );
  INV_X4 U8995 ( .A(n6674), .ZN(n6677) );
  NAND2_X2 U8996 ( .A1(n3947), .A2(n6940), .ZN(n6818) );
  NAND2_X2 U8997 ( .A1(b[20]), .A2(a[5]), .ZN(n6816) );
  INV_X4 U8998 ( .A(n6816), .ZN(n6814) );
  NAND2_X2 U8999 ( .A1(n6681), .A2(n6680), .ZN(n6684) );
  INV_X4 U9000 ( .A(n6682), .ZN(n6683) );
  AOI21_X4 U9001 ( .B1(n3967), .B2(n6684), .A(n6683), .ZN(n6879) );
  NAND2_X2 U9002 ( .A1(b[19]), .A2(a[6]), .ZN(n6810) );
  INV_X4 U9003 ( .A(n6810), .ZN(n6808) );
  NAND2_X2 U9004 ( .A1(b[18]), .A2(a[7]), .ZN(net213983) );
  NAND2_X2 U9005 ( .A1(b[17]), .A2(a[8]), .ZN(net213994) );
  INV_X4 U9006 ( .A(n6886), .ZN(n6698) );
  NAND2_X2 U9007 ( .A1(b[15]), .A2(a[10]), .ZN(n6800) );
  INV_X4 U9008 ( .A(n6800), .ZN(n6799) );
  AOI21_X4 U9009 ( .B1(n6704), .B2(n6703), .A(n6702), .ZN(n6893) );
  NAND2_X2 U9010 ( .A1(b[14]), .A2(a[11]), .ZN(n6796) );
  INV_X4 U9011 ( .A(n6796), .ZN(n6794) );
  NAND2_X2 U9012 ( .A1(b[13]), .A2(a[12]), .ZN(n6792) );
  INV_X4 U9013 ( .A(n6792), .ZN(n6790) );
  NAND2_X2 U9014 ( .A1(a[13]), .A2(b[12]), .ZN(n6784) );
  INV_X4 U9015 ( .A(n6784), .ZN(n6782) );
  INV_X4 U9016 ( .A(n6715), .ZN(n6719) );
  INV_X4 U9017 ( .A(n6716), .ZN(n6718) );
  NAND2_X2 U9018 ( .A1(a[16]), .A2(b[9]), .ZN(n6770) );
  INV_X4 U9019 ( .A(n6770), .ZN(n6765) );
  INV_X4 U9020 ( .A(n6726), .ZN(n6730) );
  INV_X4 U9021 ( .A(n6727), .ZN(n6729) );
  NAND2_X2 U9022 ( .A1(b[7]), .A2(a[18]), .ZN(n6759) );
  INV_X4 U9023 ( .A(n6759), .ZN(n6756) );
  INV_X4 U9024 ( .A(n6733), .ZN(n6737) );
  INV_X4 U9025 ( .A(n6734), .ZN(n6736) );
  OAI21_X4 U9026 ( .B1(n6737), .B2(n6736), .A(n6735), .ZN(n6912) );
  NAND2_X2 U9027 ( .A1(a[19]), .A2(b[6]), .ZN(n6754) );
  INV_X4 U9028 ( .A(n6754), .ZN(n6751) );
  INV_X4 U9029 ( .A(n6738), .ZN(n6741) );
  OAI21_X4 U9030 ( .B1(n6741), .B2(n6740), .A(n6739), .ZN(n6917) );
  NAND2_X2 U9031 ( .A1(a[20]), .A2(b[5]), .ZN(n6749) );
  INV_X4 U9032 ( .A(n6749), .ZN(n6748) );
  INV_X4 U9033 ( .A(n6742), .ZN(n6745) );
  OAI21_X4 U9034 ( .B1(n6745), .B2(n6744), .A(n6743), .ZN(net213805) );
  NAND2_X2 U9035 ( .A1(a[22]), .A2(net218538), .ZN(n6746) );
  INV_X4 U9036 ( .A(net214087), .ZN(net214089) );
  NAND2_X2 U9037 ( .A1(n6746), .A2(net214089), .ZN(net214086) );
  NAND3_X2 U9038 ( .A1(a[22]), .A2(net214087), .A3(net218534), .ZN(net213837)
         );
  NAND3_X2 U9039 ( .A1(a[21]), .A2(net214078), .A3(b[4]), .ZN(net213808) );
  NAND2_X2 U9040 ( .A1(a[21]), .A2(b[4]), .ZN(n6747) );
  INV_X4 U9041 ( .A(net214078), .ZN(net214077) );
  NAND2_X2 U9042 ( .A1(n6747), .A2(net214077), .ZN(net213806) );
  NAND2_X2 U9043 ( .A1(n6748), .A2(net214073), .ZN(n6918) );
  INV_X4 U9044 ( .A(net214073), .ZN(net214072) );
  NAND2_X2 U9045 ( .A1(n6749), .A2(net214072), .ZN(n6916) );
  NAND2_X2 U9046 ( .A1(n6918), .A2(n6916), .ZN(n6750) );
  XNOR2_X2 U9047 ( .A(n6917), .B(n6750), .ZN(n6752) );
  NAND2_X2 U9048 ( .A1(n6751), .A2(n6752), .ZN(n6913) );
  INV_X4 U9049 ( .A(n6752), .ZN(n6753) );
  NAND2_X2 U9050 ( .A1(n6913), .A2(n6911), .ZN(n6755) );
  XNOR2_X2 U9051 ( .A(n6912), .B(n6755), .ZN(n6757) );
  NAND2_X2 U9052 ( .A1(n6756), .A2(n6757), .ZN(net213850) );
  INV_X4 U9053 ( .A(n6757), .ZN(n6758) );
  NAND2_X2 U9054 ( .A1(n6759), .A2(n6758), .ZN(net213852) );
  INV_X4 U9055 ( .A(net214057), .ZN(net214059) );
  NAND2_X2 U9056 ( .A1(b[8]), .A2(a[17]), .ZN(n6760) );
  INV_X4 U9057 ( .A(n6760), .ZN(n6761) );
  NAND2_X2 U9058 ( .A1(n6761), .A2(net214057), .ZN(n6909) );
  NAND2_X2 U9059 ( .A1(n6906), .A2(n6909), .ZN(n6762) );
  XNOR2_X2 U9060 ( .A(n6763), .B(n6762), .ZN(n6764) );
  NAND2_X2 U9061 ( .A1(n6765), .A2(n6764), .ZN(n6902) );
  INV_X4 U9062 ( .A(n6766), .ZN(n6908) );
  INV_X4 U9063 ( .A(n6767), .ZN(n6907) );
  NOR2_X4 U9064 ( .A1(n6908), .A2(n6907), .ZN(n6768) );
  XNOR2_X2 U9065 ( .A(n6768), .B(n6762), .ZN(n6769) );
  NAND2_X2 U9066 ( .A1(n6770), .A2(n6769), .ZN(n6905) );
  NAND2_X2 U9067 ( .A1(n6902), .A2(n6905), .ZN(n6771) );
  XNOR2_X2 U9068 ( .A(n6772), .B(n6771), .ZN(n6775) );
  NAND2_X2 U9069 ( .A1(a[15]), .A2(b[10]), .ZN(n6774) );
  INV_X4 U9070 ( .A(n6774), .ZN(n6776) );
  NAND2_X2 U9071 ( .A1(n6776), .A2(n6775), .ZN(net213548) );
  XNOR2_X2 U9072 ( .A(net214038), .B(net214039), .ZN(n6779) );
  INV_X4 U9073 ( .A(n6779), .ZN(n6777) );
  NAND2_X2 U9074 ( .A1(a[14]), .A2(b[11]), .ZN(n6778) );
  INV_X4 U9075 ( .A(n6778), .ZN(n6780) );
  XNOR2_X2 U9076 ( .A(n6781), .B(net214033), .ZN(n6783) );
  NOR2_X4 U9077 ( .A1(net213766), .A2(net214024), .ZN(n6788) );
  NOR2_X4 U9078 ( .A1(n6789), .A2(net214022), .ZN(net213560) );
  XNOR2_X2 U9079 ( .A(n6896), .B(n6793), .ZN(n6795) );
  XNOR2_X2 U9080 ( .A(n6802), .B(n6801), .ZN(n6805) );
  NAND2_X2 U9081 ( .A1(b[16]), .A2(a[9]), .ZN(n6804) );
  INV_X4 U9082 ( .A(n6804), .ZN(n6806) );
  INV_X4 U9083 ( .A(net213995), .ZN(net213993) );
  XNOR2_X2 U9084 ( .A(n6807), .B(net213981), .ZN(n6809) );
  NAND2_X2 U9085 ( .A1(n6808), .A2(n6809), .ZN(n6881) );
  INV_X4 U9086 ( .A(n3874), .ZN(n6811) );
  XNOR2_X2 U9087 ( .A(n6813), .B(n6812), .ZN(n6815) );
  INV_X4 U9088 ( .A(n6815), .ZN(n6817) );
  XNOR2_X2 U9089 ( .A(net213969), .B(n6818), .ZN(n6820) );
  XNOR2_X2 U9090 ( .A(n6824), .B(n6823), .ZN(n6826) );
  NAND2_X2 U9091 ( .A1(b[24]), .A2(a[1]), .ZN(n6836) );
  OAI21_X4 U9092 ( .B1(n6835), .B2(n6834), .A(n6836), .ZN(n6869) );
  INV_X4 U9093 ( .A(n6836), .ZN(n6837) );
  XNOR2_X2 U9094 ( .A(n6841), .B(n6868), .ZN(n6844) );
  INV_X4 U9095 ( .A(n6844), .ZN(n6972) );
  OAI211_X2 U9096 ( .C1(n6972), .C2(n7888), .A(net218610), .B(n3405), .ZN(
        n6848) );
  AOI211_X2 U9097 ( .C1(b[25]), .C2(n6848), .A(n6847), .B(n6846), .ZN(n6867)
         );
  INV_X4 U9098 ( .A(n6852), .ZN(n6853) );
  AOI22_X2 U9099 ( .A1(n6854), .A2(n3336), .B1(a[24]), .B2(n6853), .ZN(n6990)
         );
  XNOR2_X2 U9100 ( .A(n4002), .B(b[25]), .ZN(n6991) );
  XNOR2_X2 U9101 ( .A(n6991), .B(net213919), .ZN(n6989) );
  XNOR2_X2 U9102 ( .A(n6990), .B(n6989), .ZN(n6858) );
  NAND2_X2 U9103 ( .A1(n7050), .A2(net212971), .ZN(n6857) );
  NAND2_X2 U9104 ( .A1(n7040), .A2(n6855), .ZN(n6856) );
  OAI211_X2 U9105 ( .C1(n7389), .C2(n6858), .A(n6857), .B(n6856), .ZN(n6864)
         );
  NAND2_X2 U9106 ( .A1(net218639), .A2(n6859), .ZN(n6860) );
  NOR3_X2 U9107 ( .A1(n6864), .A2(n6863), .A3(n6862), .ZN(n6865) );
  NAND3_X2 U9108 ( .A1(n6867), .A2(n6866), .A3(n6865), .ZN(result[25]) );
  INV_X4 U9109 ( .A(n6868), .ZN(n6870) );
  NAND2_X2 U9110 ( .A1(b[24]), .A2(a[2]), .ZN(n6967) );
  INV_X4 U9111 ( .A(n6967), .ZN(n6966) );
  NAND2_X2 U9112 ( .A1(a[3]), .A2(b[23]), .ZN(n6951) );
  INV_X4 U9113 ( .A(n6951), .ZN(n6950) );
  NAND2_X2 U9114 ( .A1(n6871), .A2(net213609), .ZN(n6948) );
  NAND2_X2 U9115 ( .A1(b[22]), .A2(net219055), .ZN(n6946) );
  INV_X4 U9116 ( .A(n6946), .ZN(n6944) );
  NAND3_X2 U9117 ( .A1(n6874), .A2(n6875), .A3(n6876), .ZN(net213604) );
  NAND2_X2 U9118 ( .A1(a[6]), .A2(b[20]), .ZN(net213712) );
  INV_X4 U9119 ( .A(n6877), .ZN(n6883) );
  OAI21_X4 U9120 ( .B1(n6883), .B2(n6882), .A(n6881), .ZN(net213593) );
  NAND2_X2 U9121 ( .A1(a[9]), .A2(b[17]), .ZN(n6936) );
  INV_X4 U9122 ( .A(n6936), .ZN(n6935) );
  NAND2_X2 U9123 ( .A1(a[10]), .A2(b[16]), .ZN(n6934) );
  INV_X4 U9124 ( .A(n6934), .ZN(n6933) );
  OAI21_X4 U9125 ( .B1(n6890), .B2(n6889), .A(n6888), .ZN(net213571) );
  NAND2_X2 U9126 ( .A1(a[11]), .A2(b[15]), .ZN(n6932) );
  INV_X4 U9127 ( .A(n6932), .ZN(n6931) );
  OAI21_X4 U9128 ( .B1(n6894), .B2(n6893), .A(n6892), .ZN(net213566) );
  OAI21_X4 U9129 ( .B1(n6899), .B2(n6898), .A(n3193), .ZN(net213752) );
  INV_X4 U9130 ( .A(net213867), .ZN(net213865) );
  OAI21_X4 U9131 ( .B1(net213864), .B2(net213865), .A(net213866), .ZN(
        net213547) );
  INV_X4 U9132 ( .A(n6902), .ZN(n6903) );
  AOI21_X4 U9133 ( .B1(n6905), .B2(n6904), .A(n6903), .ZN(net213541) );
  NAND2_X2 U9134 ( .A1(a[17]), .A2(b[9]), .ZN(n6929) );
  INV_X4 U9135 ( .A(n6929), .ZN(n6928) );
  OAI21_X4 U9136 ( .B1(n6908), .B2(n6907), .A(n6906), .ZN(n6910) );
  NAND2_X2 U9137 ( .A1(n6910), .A2(n6909), .ZN(net213177) );
  NAND2_X2 U9138 ( .A1(b[8]), .A2(a[18]), .ZN(n6927) );
  INV_X4 U9139 ( .A(n6927), .ZN(n6926) );
  NAND2_X2 U9140 ( .A1(b[7]), .A2(a[19]), .ZN(net213790) );
  INV_X4 U9141 ( .A(n6911), .ZN(n6915) );
  INV_X4 U9142 ( .A(n6912), .ZN(n6914) );
  OAI21_X4 U9143 ( .B1(n6915), .B2(n6914), .A(n6913), .ZN(net213533) );
  NAND2_X2 U9144 ( .A1(a[20]), .A2(b[6]), .ZN(n6925) );
  INV_X4 U9145 ( .A(n6925), .ZN(n6924) );
  INV_X4 U9146 ( .A(n6916), .ZN(n6920) );
  INV_X4 U9147 ( .A(n6917), .ZN(n6919) );
  OAI21_X4 U9148 ( .B1(n6920), .B2(n6919), .A(n6918), .ZN(net213528) );
  NAND2_X2 U9149 ( .A1(a[21]), .A2(b[5]), .ZN(n6923) );
  INV_X4 U9150 ( .A(n6923), .ZN(n6922) );
  INV_X4 U9151 ( .A(n6921), .ZN(n7219) );
  NAND2_X2 U9152 ( .A1(n7219), .A2(a[25]), .ZN(net213513) );
  NAND2_X2 U9153 ( .A1(n6922), .A2(net213802), .ZN(net213527) );
  INV_X4 U9154 ( .A(net213802), .ZN(net213801) );
  NAND2_X2 U9155 ( .A1(n6923), .A2(net213801), .ZN(net213529) );
  NAND2_X2 U9156 ( .A1(n6924), .A2(net213797), .ZN(net213532) );
  INV_X4 U9157 ( .A(net213797), .ZN(net213795) );
  NAND2_X2 U9158 ( .A1(net213795), .A2(n6925), .ZN(net213534) );
  NAND2_X2 U9159 ( .A1(n6926), .A2(net213787), .ZN(net213473) );
  INV_X4 U9160 ( .A(net213787), .ZN(net213786) );
  NAND2_X2 U9161 ( .A1(n6927), .A2(net213786), .ZN(net213178) );
  NAND2_X2 U9162 ( .A1(n6928), .A2(net213782), .ZN(net213542) );
  INV_X4 U9163 ( .A(net213782), .ZN(net213780) );
  XNOR2_X2 U9164 ( .A(net213778), .B(net213779), .ZN(net213775) );
  NAND2_X2 U9165 ( .A1(a[16]), .A2(b[10]), .ZN(net213776) );
  XNOR2_X2 U9166 ( .A(net213772), .B(net213773), .ZN(net213769) );
  NAND2_X2 U9167 ( .A1(a[15]), .A2(b[11]), .ZN(net213770) );
  INV_X4 U9168 ( .A(net213767), .ZN(net213761) );
  XNOR2_X2 U9169 ( .A(net213761), .B(net213762), .ZN(net213758) );
  NAND2_X2 U9170 ( .A1(a[14]), .A2(b[12]), .ZN(net213759) );
  NAND2_X2 U9171 ( .A1(a[12]), .A2(b[14]), .ZN(n6930) );
  NAND2_X2 U9172 ( .A1(net213745), .A2(n6931), .ZN(net213570) );
  INV_X4 U9173 ( .A(net213745), .ZN(net213743) );
  NAND2_X2 U9174 ( .A1(n6933), .A2(net213740), .ZN(net213575) );
  INV_X4 U9175 ( .A(net213740), .ZN(net213738) );
  INV_X4 U9176 ( .A(net213737), .ZN(net213734) );
  NAND2_X2 U9177 ( .A1(n6935), .A2(net213732), .ZN(net213229) );
  NAND2_X2 U9178 ( .A1(a[8]), .A2(b[18]), .ZN(net213722) );
  NAND2_X2 U9179 ( .A1(a[7]), .A2(b[19]), .ZN(n6937) );
  INV_X4 U9180 ( .A(n6937), .ZN(n6938) );
  NAND2_X2 U9181 ( .A1(n6938), .A2(net213716), .ZN(net213592) );
  INV_X4 U9182 ( .A(net213707), .ZN(net213702) );
  XNOR2_X2 U9183 ( .A(net213704), .B(net213705), .ZN(n6941) );
  XNOR2_X2 U9184 ( .A(n6943), .B(n6942), .ZN(n6945) );
  NAND2_X2 U9185 ( .A1(n6945), .A2(n6944), .ZN(net213022) );
  XNOR2_X2 U9186 ( .A(net213692), .B(n6948), .ZN(n6952) );
  INV_X4 U9187 ( .A(n6952), .ZN(n6949) );
  NAND2_X2 U9188 ( .A1(n3915), .A2(n6951), .ZN(n7011) );
  NAND2_X2 U9189 ( .A1(n7113), .A2(n7011), .ZN(n6964) );
  INV_X4 U9190 ( .A(n6953), .ZN(n6960) );
  INV_X4 U9191 ( .A(n6954), .ZN(n6959) );
  NOR2_X4 U9192 ( .A1(net213683), .A2(net213684), .ZN(n6957) );
  INV_X4 U9193 ( .A(net213680), .ZN(net213611) );
  XNOR2_X2 U9194 ( .A(n6957), .B(net213611), .ZN(n6958) );
  XNOR2_X2 U9195 ( .A(n6964), .B(n6963), .ZN(n6968) );
  XNOR2_X2 U9196 ( .A(n6969), .B(n6970), .ZN(n6971) );
  XNOR2_X2 U9197 ( .A(n6973), .B(n7105), .ZN(n6976) );
  INV_X4 U9198 ( .A(n6976), .ZN(n7029) );
  OAI211_X2 U9199 ( .C1(n7029), .C2(net218655), .A(net218608), .B(n3407), .ZN(
        n6980) );
  AOI211_X2 U9200 ( .C1(b[26]), .C2(n6980), .A(n6979), .B(n6978), .ZN(n7009)
         );
  XNOR2_X2 U9201 ( .A(n4002), .B(b[26]), .ZN(n7047) );
  INV_X4 U9202 ( .A(a[25]), .ZN(net213639) );
  OAI22_X2 U9203 ( .A1(n6991), .A2(net213639), .B1(n6990), .B2(n6989), .ZN(
        n7049) );
  XNOR2_X2 U9204 ( .A(n3337), .B(n7049), .ZN(n6998) );
  NOR2_X4 U9205 ( .A1(n6992), .A2(n3371), .ZN(n6994) );
  MUX2_X2 U9206 ( .A(net213311), .B(net213634), .S(net218556), .Z(n6993) );
  NAND2_X2 U9207 ( .A1(n6994), .A2(n6993), .ZN(n7804) );
  NAND2_X2 U9208 ( .A1(n7050), .A2(n7804), .ZN(n6997) );
  NAND2_X2 U9209 ( .A1(n7040), .A2(n6995), .ZN(n6996) );
  OAI211_X2 U9210 ( .C1(n7389), .C2(n6998), .A(n6997), .B(n6996), .ZN(n7006)
         );
  INV_X4 U9211 ( .A(n7000), .ZN(n7003) );
  NAND2_X2 U9212 ( .A1(net218639), .A2(n7001), .ZN(n7002) );
  NOR3_X2 U9213 ( .A1(n7006), .A2(n7005), .A3(n7004), .ZN(n7007) );
  NAND3_X2 U9214 ( .A1(n7009), .A2(n7008), .A3(n7007), .ZN(result[26]) );
  NAND3_X2 U9215 ( .A1(n7013), .A2(n7012), .A3(n7011), .ZN(net213251) );
  NAND2_X2 U9216 ( .A1(net219055), .A2(b[23]), .ZN(net213383) );
  NAND2_X2 U9217 ( .A1(a[9]), .A2(b[18]), .ZN(net213410) );
  NAND2_X2 U9218 ( .A1(a[26]), .A2(net218558), .ZN(n7115) );
  XNOR2_X2 U9219 ( .A(n7115), .B(n7816), .ZN(n7014) );
  INV_X4 U9220 ( .A(n7014), .ZN(n7015) );
  INV_X4 U9221 ( .A(n7017), .ZN(n7016) );
  NAND3_X4 U9222 ( .A1(n7016), .A2(a[25]), .A3(net218546), .ZN(n7125) );
  NAND2_X2 U9223 ( .A1(a[25]), .A2(net218550), .ZN(n7018) );
  NAND2_X2 U9224 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  NAND2_X2 U9225 ( .A1(n7125), .A2(n7019), .ZN(n7126) );
  XNOR2_X2 U9226 ( .A(net213152), .B(n7126), .ZN(n7020) );
  NAND3_X2 U9227 ( .A1(a[24]), .A2(n7020), .A3(net218534), .ZN(net213141) );
  NAND2_X2 U9228 ( .A1(a[24]), .A2(net218538), .ZN(n7022) );
  INV_X4 U9229 ( .A(n7020), .ZN(n7021) );
  NAND2_X2 U9230 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  XNOR2_X2 U9231 ( .A(net213380), .B(net213381), .ZN(n7024) );
  NAND2_X2 U9232 ( .A1(b[25]), .A2(a[2]), .ZN(n7107) );
  XNOR2_X2 U9233 ( .A(n3423), .B(n7107), .ZN(n7025) );
  INV_X4 U9234 ( .A(net213367), .ZN(net213364) );
  NAND3_X4 U9235 ( .A1(a[0]), .A2(b[26]), .A3(n7029), .ZN(n7101) );
  XNOR2_X2 U9236 ( .A(n7030), .B(n7101), .ZN(n7100) );
  OAI211_X2 U9237 ( .C1(n7044), .C2(n3991), .A(net218608), .B(n3406), .ZN(
        n7032) );
  NAND2_X2 U9238 ( .A1(n7033), .A2(net212010), .ZN(n7065) );
  NAND2_X2 U9239 ( .A1(net218658), .A2(net213272), .ZN(n7034) );
  NAND2_X2 U9240 ( .A1(n7034), .A2(net212094), .ZN(n7045) );
  NAND3_X2 U9241 ( .A1(n7040), .A2(a[31]), .A3(n7079), .ZN(n7037) );
  NAND2_X2 U9242 ( .A1(n7037), .A2(n7036), .ZN(net213275) );
  INV_X4 U9243 ( .A(net213275), .ZN(net212061) );
  NAND2_X2 U9244 ( .A1(n7040), .A2(n7039), .ZN(n7828) );
  INV_X4 U9245 ( .A(n7046), .ZN(n7872) );
  INV_X4 U9246 ( .A(n7047), .ZN(n7048) );
  AOI22_X2 U9247 ( .A1(n7049), .A2(n3337), .B1(a[26]), .B2(n7048), .ZN(n7093)
         );
  XNOR2_X2 U9248 ( .A(n4002), .B(b[27]), .ZN(n7095) );
  XNOR2_X2 U9249 ( .A(n7095), .B(n7054), .ZN(n7092) );
  XNOR2_X2 U9250 ( .A(n7093), .B(n7092), .ZN(n7052) );
  NAND2_X2 U9251 ( .A1(n7050), .A2(net212007), .ZN(n7051) );
  OAI221_X2 U9252 ( .B1(n7872), .B2(n7053), .C1(n7389), .C2(n7052), .A(n7051), 
        .ZN(n7062) );
  INV_X4 U9253 ( .A(n7055), .ZN(n7056) );
  NAND2_X2 U9254 ( .A1(net218639), .A2(n7056), .ZN(n7057) );
  NOR3_X2 U9255 ( .A1(n7062), .A2(n7061), .A3(n7060), .ZN(n7063) );
  NAND4_X2 U9256 ( .A1(n7066), .A2(n7065), .A3(n7064), .A4(n7063), .ZN(
        result[27]) );
  MUX2_X2 U9257 ( .A(n7816), .B(net213311), .S(net218556), .Z(n7071) );
  INV_X4 U9258 ( .A(n7068), .ZN(n7069) );
  INV_X4 U9259 ( .A(n7072), .ZN(n7088) );
  INV_X4 U9260 ( .A(n7073), .ZN(n7075) );
  OAI22_X2 U9261 ( .A1(n3993), .A2(n7075), .B1(n7074), .B2(n7869), .ZN(n7076)
         );
  MUX2_X2 U9262 ( .A(n7086), .B(n7085), .S(b[4]), .Z(n7087) );
  NAND2_X2 U9263 ( .A1(n7088), .A2(n7087), .ZN(n7091) );
  OAI22_X2 U9264 ( .A1(n7206), .A2(net218610), .B1(n7089), .B2(net218640), 
        .ZN(n7090) );
  XNOR2_X2 U9265 ( .A(n4002), .B(b[28]), .ZN(n7383) );
  XNOR2_X2 U9266 ( .A(n7383), .B(n7206), .ZN(n7382) );
  INV_X4 U9267 ( .A(a[27]), .ZN(n7094) );
  OAI22_X2 U9268 ( .A1(n7095), .A2(n7094), .B1(n7093), .B2(n7092), .ZN(n7386)
         );
  XNOR2_X2 U9269 ( .A(n7382), .B(n7386), .ZN(n7096) );
  NAND2_X2 U9270 ( .A1(n7096), .A2(n3990), .ZN(n7213) );
  NAND2_X2 U9271 ( .A1(n7866), .A2(n7097), .ZN(n7379) );
  NAND2_X2 U9272 ( .A1(n7828), .A2(n7379), .ZN(n7098) );
  NOR3_X4 U9273 ( .A1(n7100), .A2(net213272), .A3(net218496), .ZN(net212697)
         );
  INV_X4 U9274 ( .A(n7101), .ZN(n7103) );
  NAND2_X2 U9275 ( .A1(net212704), .A2(n3191), .ZN(n7205) );
  NAND2_X2 U9276 ( .A1(b[26]), .A2(a[2]), .ZN(n7202) );
  INV_X4 U9277 ( .A(n7202), .ZN(n7200) );
  XNOR2_X2 U9278 ( .A(n7108), .B(n7107), .ZN(n7106) );
  XNOR2_X2 U9279 ( .A(n7106), .B(net219657), .ZN(n7236) );
  INV_X4 U9280 ( .A(n7107), .ZN(n7110) );
  INV_X4 U9281 ( .A(n7233), .ZN(n7237) );
  NAND2_X2 U9282 ( .A1(b[25]), .A2(a[3]), .ZN(n7197) );
  INV_X4 U9283 ( .A(n7197), .ZN(n7195) );
  NAND2_X2 U9284 ( .A1(b[24]), .A2(net219055), .ZN(n7192) );
  NAND2_X2 U9285 ( .A1(a[11]), .A2(b[17]), .ZN(n7189) );
  INV_X4 U9286 ( .A(n7189), .ZN(n7187) );
  INV_X4 U9287 ( .A(net213070), .ZN(net213072) );
  XNOR2_X2 U9288 ( .A(net212906), .B(n7246), .ZN(n7174) );
  NAND2_X2 U9289 ( .A1(net212900), .A2(net220199), .ZN(n7167) );
  NAND2_X2 U9290 ( .A1(a[19]), .A2(b[9]), .ZN(n7155) );
  INV_X4 U9291 ( .A(n7155), .ZN(n7153) );
  NAND2_X2 U9292 ( .A1(b[8]), .A2(a[20]), .ZN(n7151) );
  INV_X4 U9293 ( .A(n7151), .ZN(n7148) );
  NAND2_X2 U9294 ( .A1(b[7]), .A2(a[21]), .ZN(n7146) );
  INV_X4 U9295 ( .A(n7146), .ZN(n7143) );
  INV_X4 U9296 ( .A(n7140), .ZN(n7137) );
  NAND2_X2 U9297 ( .A1(a[24]), .A2(b[4]), .ZN(n7133) );
  NAND2_X2 U9298 ( .A1(a[25]), .A2(net218538), .ZN(n7129) );
  NAND2_X2 U9299 ( .A1(a[26]), .A2(net218550), .ZN(n7122) );
  OAI21_X4 U9300 ( .B1(n7115), .B2(n7816), .A(n7114), .ZN(n7116) );
  INV_X4 U9301 ( .A(n7864), .ZN(n7117) );
  NAND2_X2 U9302 ( .A1(n7117), .A2(a[27]), .ZN(n7271) );
  NAND2_X2 U9303 ( .A1(a[27]), .A2(net218556), .ZN(n7118) );
  NAND2_X2 U9304 ( .A1(n7118), .A2(n7217), .ZN(n7119) );
  NAND2_X2 U9305 ( .A1(n7271), .A2(n7119), .ZN(n7272) );
  INV_X4 U9306 ( .A(n7272), .ZN(n7120) );
  XNOR2_X2 U9307 ( .A(n7273), .B(n7120), .ZN(n7123) );
  INV_X4 U9308 ( .A(n7123), .ZN(n7121) );
  NAND2_X2 U9309 ( .A1(n7122), .A2(n7121), .ZN(n7124) );
  NAND3_X2 U9310 ( .A1(a[26]), .A2(n7123), .A3(net218546), .ZN(n7268) );
  NAND2_X2 U9311 ( .A1(n7124), .A2(n7268), .ZN(n7269) );
  INV_X4 U9312 ( .A(net213152), .ZN(net213149) );
  NAND2_X2 U9313 ( .A1(n7129), .A2(n7128), .ZN(n7131) );
  NAND3_X2 U9314 ( .A1(a[25]), .A2(n7130), .A3(net218534), .ZN(n7266) );
  INV_X4 U9315 ( .A(net213138), .ZN(net212871) );
  INV_X4 U9316 ( .A(n7134), .ZN(n7132) );
  NAND2_X2 U9317 ( .A1(n7133), .A2(n7132), .ZN(n7135) );
  NAND3_X2 U9318 ( .A1(a[24]), .A2(n7134), .A3(b[4]), .ZN(n7264) );
  INV_X4 U9319 ( .A(net213127), .ZN(net212874) );
  XNOR2_X2 U9320 ( .A(n7136), .B(net212874), .ZN(n7138) );
  NAND2_X2 U9321 ( .A1(n7137), .A2(n7138), .ZN(n7292) );
  INV_X4 U9322 ( .A(n7138), .ZN(n7139) );
  XNOR2_X2 U9323 ( .A(net212842), .B(n7141), .ZN(n7142) );
  INV_X4 U9324 ( .A(net213111), .ZN(net212877) );
  NAND2_X2 U9325 ( .A1(n7143), .A2(n7144), .ZN(n7300) );
  INV_X4 U9326 ( .A(n7144), .ZN(n7145) );
  XNOR2_X2 U9327 ( .A(net212826), .B(n7147), .ZN(n7149) );
  NAND2_X2 U9328 ( .A1(n7148), .A2(n7149), .ZN(n7260) );
  INV_X4 U9329 ( .A(n7149), .ZN(n7150) );
  NAND2_X2 U9330 ( .A1(n7151), .A2(n7150), .ZN(n7259) );
  NAND2_X2 U9331 ( .A1(n7153), .A2(n7154), .ZN(n7257) );
  NAND2_X2 U9332 ( .A1(n3772), .A2(n7155), .ZN(n7256) );
  XNOR2_X2 U9333 ( .A(net212888), .B(n7156), .ZN(n7159) );
  INV_X4 U9334 ( .A(n7159), .ZN(n7157) );
  NAND2_X2 U9335 ( .A1(a[18]), .A2(b[10]), .ZN(n7158) );
  INV_X4 U9336 ( .A(n7158), .ZN(n7160) );
  NAND2_X2 U9337 ( .A1(n7160), .A2(n7159), .ZN(n7254) );
  XNOR2_X2 U9338 ( .A(net212893), .B(n7161), .ZN(n7164) );
  INV_X4 U9339 ( .A(n7164), .ZN(n7162) );
  NAND2_X2 U9340 ( .A1(a[17]), .A2(b[11]), .ZN(n7163) );
  INV_X4 U9341 ( .A(n7163), .ZN(n7165) );
  NAND2_X2 U9342 ( .A1(n7165), .A2(n7164), .ZN(n7249) );
  XNOR2_X2 U9343 ( .A(n7167), .B(n7166), .ZN(n7168) );
  OAI21_X4 U9344 ( .B1(n3328), .B2(n3957), .A(net212636), .ZN(n7396) );
  XNOR2_X2 U9345 ( .A(net212634), .B(n7396), .ZN(n7171) );
  NAND2_X2 U9346 ( .A1(b[13]), .A2(a[15]), .ZN(n7170) );
  NAND2_X2 U9347 ( .A1(n7169), .A2(n7170), .ZN(n7248) );
  INV_X4 U9348 ( .A(n7170), .ZN(n7172) );
  NAND2_X2 U9349 ( .A1(n7248), .A2(n7500), .ZN(n7244) );
  INV_X4 U9350 ( .A(n7244), .ZN(n7173) );
  XNOR2_X2 U9351 ( .A(n3779), .B(n7173), .ZN(n7175) );
  NAND2_X2 U9352 ( .A1(a[13]), .A2(b[15]), .ZN(n7178) );
  INV_X4 U9353 ( .A(n7178), .ZN(n7176) );
  NAND3_X2 U9354 ( .A1(n7177), .A2(n7245), .A3(n7176), .ZN(n7242) );
  INV_X4 U9355 ( .A(n7177), .ZN(n7179) );
  OAI21_X4 U9356 ( .B1(n7179), .B2(n7180), .A(n7178), .ZN(n7241) );
  NAND2_X2 U9357 ( .A1(n7242), .A2(n7241), .ZN(n7181) );
  XNOR2_X2 U9358 ( .A(net212911), .B(n7181), .ZN(n7184) );
  NAND2_X2 U9359 ( .A1(a[12]), .A2(b[16]), .ZN(n7183) );
  INV_X4 U9360 ( .A(n7183), .ZN(n7185) );
  NAND2_X2 U9361 ( .A1(n7185), .A2(n7184), .ZN(n7239) );
  XNOR2_X2 U9362 ( .A(net212916), .B(n7186), .ZN(n7188) );
  NAND2_X2 U9363 ( .A1(n7187), .A2(n7188), .ZN(net212920) );
  INV_X4 U9364 ( .A(n7188), .ZN(n7190) );
  XNOR2_X2 U9365 ( .A(net213012), .B(n3476), .ZN(n7193) );
  INV_X4 U9366 ( .A(n7193), .ZN(n7191) );
  INV_X4 U9367 ( .A(n7192), .ZN(n7194) );
  XNOR2_X2 U9368 ( .A(net213005), .B(net213006), .ZN(n7196) );
  NAND2_X2 U9369 ( .A1(n3768), .A2(n7195), .ZN(net212443) );
  INV_X4 U9370 ( .A(n7196), .ZN(n7198) );
  INV_X4 U9371 ( .A(net213000), .ZN(net212999) );
  XNOR2_X2 U9372 ( .A(n7199), .B(net212999), .ZN(n7201) );
  NAND2_X2 U9373 ( .A1(n7200), .A2(n7201), .ZN(net212700) );
  INV_X4 U9374 ( .A(n7201), .ZN(n7203) );
  XNOR2_X2 U9375 ( .A(n7205), .B(n7204), .ZN(net212696) );
  XNOR2_X2 U9376 ( .A(net212991), .B(net212697), .ZN(n7375) );
  NAND2_X2 U9377 ( .A1(net218658), .A2(net212989), .ZN(n7208) );
  NAND4_X2 U9378 ( .A1(n7211), .A2(n7213), .A3(n7212), .A4(n7214), .ZN(
        result[28]) );
  NAND2_X2 U9379 ( .A1(n7216), .A2(n7215), .ZN(n7220) );
  INV_X4 U9380 ( .A(net212971), .ZN(net212970) );
  INV_X4 U9381 ( .A(n7222), .ZN(n7223) );
  MUX2_X2 U9382 ( .A(n7227), .B(n3379), .S(b[4]), .Z(n7228) );
  NAND2_X2 U9383 ( .A1(b[22]), .A2(a[7]), .ZN(net212738) );
  INV_X4 U9384 ( .A(net212738), .ZN(net212740) );
  INV_X4 U9385 ( .A(net220079), .ZN(net212741) );
  NAND2_X2 U9386 ( .A1(a[8]), .A2(b[21]), .ZN(n7372) );
  INV_X4 U9387 ( .A(n7372), .ZN(n7371) );
  NAND2_X2 U9388 ( .A1(a[9]), .A2(b[20]), .ZN(n7369) );
  INV_X4 U9389 ( .A(n7369), .ZN(n7368) );
  OAI21_X4 U9390 ( .B1(net212927), .B2(net212928), .A(net219674), .ZN(n7542)
         );
  NAND2_X2 U9391 ( .A1(a[10]), .A2(b[19]), .ZN(n7366) );
  INV_X4 U9392 ( .A(n7366), .ZN(n7364) );
  NAND2_X2 U9393 ( .A1(a[11]), .A2(b[18]), .ZN(n7361) );
  INV_X4 U9394 ( .A(n7361), .ZN(n7359) );
  NAND2_X2 U9395 ( .A1(a[12]), .A2(b[17]), .ZN(n7356) );
  INV_X4 U9396 ( .A(n7356), .ZN(n7354) );
  INV_X4 U9397 ( .A(n7238), .ZN(n7240) );
  INV_X4 U9398 ( .A(net212916), .ZN(net212914) );
  OAI21_X4 U9399 ( .B1(n7240), .B2(net212914), .A(n3929), .ZN(n7526) );
  NAND2_X2 U9400 ( .A1(a[13]), .A2(b[16]), .ZN(n7351) );
  INV_X4 U9401 ( .A(n7351), .ZN(n7349) );
  OAI21_X4 U9402 ( .B1(n7243), .B2(net212909), .A(n7242), .ZN(n7517) );
  XNOR2_X2 U9403 ( .A(net212906), .B(n7244), .ZN(n7247) );
  OAI21_X4 U9404 ( .B1(n7247), .B2(n7246), .A(n7245), .ZN(n7512) );
  NAND2_X2 U9405 ( .A1(a[15]), .A2(b[14]), .ZN(n7339) );
  INV_X4 U9406 ( .A(n7339), .ZN(n7337) );
  NAND2_X2 U9407 ( .A1(n7501), .A2(n7500), .ZN(n7336) );
  NAND2_X2 U9408 ( .A1(b[13]), .A2(a[16]), .ZN(n7333) );
  INV_X4 U9409 ( .A(n7333), .ZN(n7332) );
  NAND2_X2 U9410 ( .A1(net220199), .A2(net212900), .ZN(n7251) );
  AOI21_X4 U9411 ( .B1(n7252), .B2(n7251), .A(n7250), .ZN(n7492) );
  INV_X4 U9412 ( .A(n7492), .ZN(n7323) );
  NAND2_X2 U9413 ( .A1(a[18]), .A2(b[11]), .ZN(n7320) );
  INV_X4 U9414 ( .A(n7320), .ZN(n7318) );
  INV_X4 U9415 ( .A(n7253), .ZN(n7255) );
  INV_X4 U9416 ( .A(net212893), .ZN(net212891) );
  NAND2_X2 U9417 ( .A1(a[19]), .A2(b[10]), .ZN(n7316) );
  INV_X4 U9418 ( .A(n7316), .ZN(n7314) );
  INV_X4 U9419 ( .A(n7256), .ZN(n7258) );
  INV_X4 U9420 ( .A(net212888), .ZN(net212886) );
  NAND2_X2 U9421 ( .A1(a[20]), .A2(b[9]), .ZN(n7311) );
  INV_X4 U9422 ( .A(n7311), .ZN(n7309) );
  INV_X4 U9423 ( .A(n7259), .ZN(n7261) );
  NAND2_X2 U9424 ( .A1(b[8]), .A2(a[21]), .ZN(n7307) );
  INV_X4 U9425 ( .A(n7307), .ZN(n7304) );
  OAI21_X4 U9426 ( .B1(net212877), .B2(n7263), .A(n7262), .ZN(n7416) );
  NAND2_X2 U9427 ( .A1(a[23]), .A2(b[6]), .ZN(n7296) );
  INV_X4 U9428 ( .A(n7296), .ZN(n7294) );
  OAI21_X4 U9429 ( .B1(net212874), .B2(n7265), .A(n3887), .ZN(n7455) );
  NAND2_X2 U9430 ( .A1(a[25]), .A2(b[4]), .ZN(n7287) );
  NAND2_X2 U9431 ( .A1(a[28]), .A2(net218558), .ZN(n7434) );
  XNOR2_X2 U9432 ( .A(n7434), .B(n7817), .ZN(n7274) );
  INV_X4 U9433 ( .A(n7274), .ZN(n7276) );
  OAI21_X4 U9434 ( .B1(n7273), .B2(n7272), .A(n7271), .ZN(n7275) );
  NAND2_X2 U9435 ( .A1(n7276), .A2(n7275), .ZN(n7433) );
  OAI21_X4 U9436 ( .B1(n7276), .B2(n7275), .A(n7433), .ZN(n7278) );
  INV_X4 U9437 ( .A(n7278), .ZN(n7277) );
  NAND3_X4 U9438 ( .A1(n7277), .A2(a[27]), .A3(net218546), .ZN(n7430) );
  NAND2_X2 U9439 ( .A1(a[27]), .A2(net218550), .ZN(n7279) );
  NAND2_X2 U9440 ( .A1(n7279), .A2(n7278), .ZN(n7428) );
  NAND2_X2 U9441 ( .A1(n7430), .A2(n7428), .ZN(n7280) );
  XNOR2_X2 U9442 ( .A(n7429), .B(n7280), .ZN(n7283) );
  INV_X4 U9443 ( .A(n7283), .ZN(n7281) );
  NAND2_X2 U9444 ( .A1(a[26]), .A2(net218540), .ZN(n7282) );
  NAND2_X2 U9445 ( .A1(n7281), .A2(n7282), .ZN(n7423) );
  INV_X4 U9446 ( .A(n7282), .ZN(n7284) );
  NAND2_X2 U9447 ( .A1(n7284), .A2(n7283), .ZN(n7425) );
  NAND2_X2 U9448 ( .A1(n7423), .A2(n7425), .ZN(n7285) );
  XNOR2_X2 U9449 ( .A(n7424), .B(n7285), .ZN(n7288) );
  INV_X4 U9450 ( .A(n7288), .ZN(n7286) );
  NAND2_X2 U9451 ( .A1(n7287), .A2(n7286), .ZN(n7289) );
  NAND3_X2 U9452 ( .A1(a[25]), .A2(n7288), .A3(b[4]), .ZN(n7456) );
  XNOR2_X2 U9453 ( .A(n7455), .B(n7457), .ZN(n7290) );
  OAI21_X4 U9454 ( .B1(n3948), .B2(n3324), .A(n7420), .ZN(n7421) );
  INV_X4 U9455 ( .A(net212842), .ZN(net212840) );
  OAI21_X4 U9456 ( .B1(n3760), .B2(net212840), .A(n7292), .ZN(n7293) );
  INV_X4 U9457 ( .A(n7293), .ZN(n7422) );
  NAND2_X2 U9458 ( .A1(n7294), .A2(n7295), .ZN(n7417) );
  NAND2_X2 U9459 ( .A1(n3925), .A2(n7296), .ZN(n7415) );
  XNOR2_X2 U9460 ( .A(n7416), .B(n7297), .ZN(n7298) );
  OAI21_X4 U9461 ( .B1(n3323), .B2(n3876), .A(n7412), .ZN(n7413) );
  INV_X4 U9462 ( .A(n7299), .ZN(n7301) );
  INV_X4 U9463 ( .A(net212826), .ZN(net212824) );
  OAI21_X4 U9464 ( .B1(n7301), .B2(net212824), .A(n7300), .ZN(n7302) );
  INV_X4 U9465 ( .A(n7302), .ZN(n7414) );
  XNOR2_X2 U9466 ( .A(n7303), .B(n7414), .ZN(n7305) );
  NAND2_X2 U9467 ( .A1(n7304), .A2(n7305), .ZN(n7409) );
  INV_X4 U9468 ( .A(n7305), .ZN(n7306) );
  NAND2_X2 U9469 ( .A1(n7307), .A2(n7306), .ZN(n7407) );
  NAND2_X2 U9470 ( .A1(n7409), .A2(n7407), .ZN(n7308) );
  XNOR2_X2 U9471 ( .A(n7408), .B(n7308), .ZN(n7310) );
  NAND2_X2 U9472 ( .A1(n7309), .A2(n7310), .ZN(n7484) );
  INV_X4 U9473 ( .A(n7310), .ZN(n7312) );
  NAND2_X2 U9474 ( .A1(n7316), .A2(n3933), .ZN(n7401) );
  XNOR2_X2 U9475 ( .A(n7402), .B(n7317), .ZN(n7319) );
  NAND2_X2 U9476 ( .A1(n7318), .A2(n7319), .ZN(n7491) );
  INV_X4 U9477 ( .A(n7319), .ZN(n7321) );
  NAND2_X2 U9478 ( .A1(n7321), .A2(n7320), .ZN(n7490) );
  XNOR2_X2 U9479 ( .A(n7323), .B(n7322), .ZN(n7326) );
  INV_X4 U9480 ( .A(n7326), .ZN(n7324) );
  NAND2_X2 U9481 ( .A1(a[17]), .A2(b[12]), .ZN(n7325) );
  INV_X4 U9482 ( .A(n7325), .ZN(n7327) );
  NAND2_X2 U9483 ( .A1(n7327), .A2(n3901), .ZN(n7398) );
  NAND2_X2 U9484 ( .A1(n7395), .A2(n7398), .ZN(n7330) );
  NAND2_X2 U9485 ( .A1(n7396), .A2(net212636), .ZN(n7328) );
  XNOR2_X2 U9486 ( .A(n7330), .B(n7329), .ZN(n7334) );
  INV_X4 U9487 ( .A(n7334), .ZN(n7331) );
  NAND2_X2 U9488 ( .A1(n7334), .A2(n7333), .ZN(n7502) );
  XNOR2_X2 U9489 ( .A(n7336), .B(n7335), .ZN(n7338) );
  NAND2_X2 U9490 ( .A1(n7514), .A2(n7513), .ZN(n7341) );
  XNOR2_X2 U9491 ( .A(n7342), .B(n7341), .ZN(n7343) );
  NAND2_X2 U9492 ( .A1(a[14]), .A2(b[15]), .ZN(n7344) );
  INV_X4 U9493 ( .A(n7344), .ZN(n7347) );
  NAND2_X2 U9494 ( .A1(n7513), .A2(n7514), .ZN(n7345) );
  XNOR2_X2 U9495 ( .A(n7345), .B(n7512), .ZN(n7346) );
  XNOR2_X2 U9496 ( .A(n7517), .B(n7348), .ZN(n7350) );
  NAND2_X2 U9497 ( .A1(n7349), .A2(n7350), .ZN(n7527) );
  INV_X4 U9498 ( .A(n7350), .ZN(n7352) );
  XNOR2_X2 U9499 ( .A(n7526), .B(n7353), .ZN(n7355) );
  NAND2_X2 U9500 ( .A1(n7354), .A2(n7355), .ZN(n7531) );
  INV_X4 U9501 ( .A(n7355), .ZN(n7357) );
  XNOR2_X2 U9502 ( .A(net212495), .B(n7358), .ZN(n7360) );
  NAND2_X2 U9503 ( .A1(n7359), .A2(n7360), .ZN(n7539) );
  INV_X4 U9504 ( .A(n7360), .ZN(n7362) );
  XNOR2_X2 U9505 ( .A(net212485), .B(n7363), .ZN(n7365) );
  NAND2_X2 U9506 ( .A1(n7371), .A2(n3913), .ZN(n7554) );
  INV_X4 U9507 ( .A(n3913), .ZN(n7373) );
  XNOR2_X2 U9508 ( .A(net212741), .B(n7374), .ZN(net212739) );
  NAND2_X2 U9509 ( .A1(net212693), .A2(net212694), .ZN(net212686) );
  INV_X4 U9510 ( .A(net212686), .ZN(net212689) );
  INV_X4 U9511 ( .A(net212694), .ZN(net212691) );
  INV_X4 U9512 ( .A(net212685), .ZN(net212690) );
  OAI21_X4 U9513 ( .B1(net212690), .B2(net212689), .A(net212688), .ZN(
        net212411) );
  NOR2_X4 U9514 ( .A1(net218614), .A2(n7376), .ZN(net212681) );
  NOR2_X4 U9515 ( .A1(n7387), .A2(net218608), .ZN(n7377) );
  AOI21_X4 U9516 ( .B1(net212679), .B2(b[29]), .A(n7377), .ZN(n7393) );
  INV_X4 U9517 ( .A(n7379), .ZN(n7856) );
  NAND2_X2 U9518 ( .A1(n7856), .A2(n7380), .ZN(net212674) );
  INV_X4 U9519 ( .A(n7382), .ZN(n7385) );
  INV_X4 U9520 ( .A(n7383), .ZN(n7384) );
  AOI22_X2 U9521 ( .A1(n7386), .A2(n7385), .B1(a[28]), .B2(n7384), .ZN(n7841)
         );
  XNOR2_X2 U9522 ( .A(n4002), .B(b[29]), .ZN(n7843) );
  XNOR2_X2 U9523 ( .A(n7843), .B(n7387), .ZN(n7840) );
  XNOR2_X2 U9524 ( .A(n7841), .B(n7840), .ZN(n7388) );
  NAND3_X2 U9525 ( .A1(n7394), .A2(n7393), .A3(n7392), .ZN(n7897) );
  NAND2_X2 U9526 ( .A1(b[25]), .A2(a[5]), .ZN(n7571) );
  XNOR2_X2 U9527 ( .A(net212134), .B(n7571), .ZN(n7565) );
  INV_X4 U9528 ( .A(n7395), .ZN(n7400) );
  AOI21_X4 U9529 ( .B1(n7397), .B2(net212634), .A(net212635), .ZN(n7399) );
  OAI21_X4 U9530 ( .B1(n7400), .B2(n7399), .A(n7398), .ZN(n7598) );
  INV_X4 U9531 ( .A(n7598), .ZN(n7594) );
  NAND2_X2 U9532 ( .A1(b[13]), .A2(a[17]), .ZN(n7593) );
  XNOR2_X2 U9533 ( .A(n7594), .B(n7593), .ZN(n7499) );
  INV_X4 U9534 ( .A(n7401), .ZN(n7405) );
  INV_X4 U9535 ( .A(n7402), .ZN(n7404) );
  OAI21_X4 U9536 ( .B1(n7405), .B2(n7404), .A(n7403), .ZN(n7406) );
  INV_X4 U9537 ( .A(n7406), .ZN(n7730) );
  NAND2_X2 U9538 ( .A1(a[19]), .A2(b[11]), .ZN(n7600) );
  XNOR2_X2 U9539 ( .A(n7730), .B(n7600), .ZN(n7489) );
  INV_X4 U9540 ( .A(n7407), .ZN(n7411) );
  INV_X4 U9541 ( .A(n7408), .ZN(n7410) );
  OAI21_X4 U9542 ( .B1(n7411), .B2(n7410), .A(n7409), .ZN(n7476) );
  OAI21_X4 U9543 ( .B1(n7414), .B2(n7413), .A(n7412), .ZN(n7618) );
  NAND2_X2 U9544 ( .A1(a[23]), .A2(b[7]), .ZN(n7473) );
  INV_X4 U9545 ( .A(n7473), .ZN(n7470) );
  INV_X4 U9546 ( .A(n7415), .ZN(n7419) );
  INV_X4 U9547 ( .A(n7416), .ZN(n7418) );
  OAI21_X4 U9548 ( .B1(n7422), .B2(n7421), .A(n7420), .ZN(n7623) );
  NAND2_X2 U9549 ( .A1(a[26]), .A2(b[4]), .ZN(n7454) );
  INV_X4 U9550 ( .A(n7454), .ZN(n7451) );
  INV_X4 U9551 ( .A(n7423), .ZN(n7427) );
  INV_X4 U9552 ( .A(n7424), .ZN(n7426) );
  OAI21_X4 U9553 ( .B1(n7427), .B2(n7426), .A(n7425), .ZN(n7631) );
  INV_X4 U9554 ( .A(n7428), .ZN(n7432) );
  INV_X4 U9555 ( .A(n7429), .ZN(n7431) );
  OAI21_X4 U9556 ( .B1(n7432), .B2(n7431), .A(n7430), .ZN(n7633) );
  NAND2_X2 U9557 ( .A1(a[28]), .A2(net218550), .ZN(n7444) );
  INV_X4 U9558 ( .A(n7444), .ZN(n7441) );
  INV_X4 U9559 ( .A(n7637), .ZN(n7440) );
  NAND2_X2 U9560 ( .A1(a[29]), .A2(net218556), .ZN(n7439) );
  INV_X4 U9561 ( .A(n7439), .ZN(n7435) );
  NAND2_X2 U9562 ( .A1(n7436), .A2(n7435), .ZN(n7695) );
  INV_X4 U9563 ( .A(n7695), .ZN(n7437) );
  AOI21_X4 U9564 ( .B1(n7439), .B2(n7438), .A(n7437), .ZN(n7638) );
  XNOR2_X2 U9565 ( .A(n7440), .B(n7638), .ZN(n7442) );
  NAND2_X2 U9566 ( .A1(n7441), .A2(n7442), .ZN(n7634) );
  INV_X4 U9567 ( .A(n7442), .ZN(n7443) );
  NAND2_X2 U9568 ( .A1(n7444), .A2(n7443), .ZN(n7632) );
  NAND2_X2 U9569 ( .A1(n7634), .A2(n7632), .ZN(n7445) );
  XNOR2_X2 U9570 ( .A(n7633), .B(n7445), .ZN(n7448) );
  INV_X4 U9571 ( .A(n7448), .ZN(n7446) );
  NAND2_X2 U9572 ( .A1(a[27]), .A2(net218540), .ZN(n7447) );
  NAND2_X2 U9573 ( .A1(n7446), .A2(n7447), .ZN(n7630) );
  INV_X4 U9574 ( .A(n7447), .ZN(n7449) );
  NAND2_X2 U9575 ( .A1(n7449), .A2(n7448), .ZN(n7628) );
  NAND2_X2 U9576 ( .A1(n7630), .A2(n7628), .ZN(n7450) );
  XNOR2_X2 U9577 ( .A(n7631), .B(n7450), .ZN(n7452) );
  NAND2_X2 U9578 ( .A1(n7451), .A2(n7452), .ZN(n7627) );
  INV_X4 U9579 ( .A(n7452), .ZN(n7453) );
  NAND2_X2 U9580 ( .A1(n7454), .A2(n7453), .ZN(n7459) );
  INV_X4 U9581 ( .A(n7455), .ZN(n7458) );
  NAND3_X2 U9582 ( .A1(n7460), .A2(n7627), .A3(n7459), .ZN(n7711) );
  INV_X4 U9583 ( .A(n7463), .ZN(n7462) );
  NAND2_X2 U9584 ( .A1(a[25]), .A2(b[5]), .ZN(n7464) );
  INV_X4 U9585 ( .A(n7464), .ZN(n7461) );
  NAND2_X2 U9586 ( .A1(n7462), .A2(n7461), .ZN(n7624) );
  NAND2_X2 U9587 ( .A1(n7464), .A2(n7463), .ZN(n7622) );
  NAND2_X2 U9588 ( .A1(n7624), .A2(n7622), .ZN(n7465) );
  XNOR2_X2 U9589 ( .A(n7623), .B(n7465), .ZN(n7619) );
  NAND2_X2 U9590 ( .A1(a[24]), .A2(b[6]), .ZN(n7620) );
  XNOR2_X2 U9591 ( .A(n7619), .B(n7620), .ZN(n7467) );
  NAND2_X2 U9592 ( .A1(n7466), .A2(n7467), .ZN(n7471) );
  INV_X4 U9593 ( .A(n7466), .ZN(n7469) );
  INV_X4 U9594 ( .A(n7467), .ZN(n7468) );
  NAND2_X2 U9595 ( .A1(n7469), .A2(n7468), .ZN(n7472) );
  NAND3_X2 U9596 ( .A1(n7470), .A2(n7471), .A3(n7472), .ZN(n7615) );
  INV_X4 U9597 ( .A(n7471), .ZN(n7718) );
  INV_X4 U9598 ( .A(n7472), .ZN(n7474) );
  OAI21_X4 U9599 ( .B1(n7718), .B2(n7474), .A(n7473), .ZN(n7617) );
  NAND2_X2 U9600 ( .A1(n7615), .A2(n7617), .ZN(n7475) );
  XNOR2_X2 U9601 ( .A(n7618), .B(n7475), .ZN(n7612) );
  NAND2_X2 U9602 ( .A1(a[22]), .A2(b[8]), .ZN(n7613) );
  XNOR2_X2 U9603 ( .A(n7612), .B(n7613), .ZN(n7477) );
  NAND2_X2 U9604 ( .A1(n7476), .A2(n7477), .ZN(n7723) );
  INV_X4 U9605 ( .A(n7476), .ZN(n7479) );
  INV_X4 U9606 ( .A(n7477), .ZN(n7478) );
  NAND2_X2 U9607 ( .A1(n7479), .A2(n7478), .ZN(n7480) );
  NAND4_X2 U9608 ( .A1(a[21]), .A2(n7723), .A3(b[9]), .A4(n7480), .ZN(n7609)
         );
  INV_X4 U9609 ( .A(n7609), .ZN(n7481) );
  AOI22_X2 U9610 ( .A1(n7723), .A2(n7480), .B1(a[21]), .B2(b[9]), .ZN(n7611)
         );
  NOR2_X4 U9611 ( .A1(n7481), .A2(n7611), .ZN(n7488) );
  INV_X4 U9612 ( .A(n7482), .ZN(n7486) );
  INV_X4 U9613 ( .A(n7483), .ZN(n7485) );
  INV_X4 U9614 ( .A(n7487), .ZN(n7610) );
  XNOR2_X2 U9615 ( .A(n7488), .B(n7610), .ZN(n7606) );
  NAND2_X2 U9616 ( .A1(a[20]), .A2(b[10]), .ZN(n7607) );
  XNOR2_X2 U9617 ( .A(n7606), .B(n7607), .ZN(n7601) );
  INV_X4 U9618 ( .A(n7601), .ZN(n7729) );
  XNOR2_X2 U9619 ( .A(n7489), .B(n7729), .ZN(n7494) );
  INV_X4 U9620 ( .A(n7494), .ZN(n7497) );
  INV_X4 U9621 ( .A(n7494), .ZN(n7495) );
  NAND2_X2 U9622 ( .A1(n7495), .A2(n7496), .ZN(n7604) );
  OAI21_X4 U9623 ( .B1(n7497), .B2(n7496), .A(n7604), .ZN(n7736) );
  NAND2_X2 U9624 ( .A1(a[18]), .A2(b[12]), .ZN(n7735) );
  XNOR2_X2 U9625 ( .A(n7736), .B(n7735), .ZN(n7498) );
  INV_X4 U9626 ( .A(n7498), .ZN(n7599) );
  XNOR2_X2 U9627 ( .A(n7499), .B(n7599), .ZN(n7508) );
  INV_X4 U9628 ( .A(n7500), .ZN(n7504) );
  INV_X4 U9629 ( .A(n7501), .ZN(n7503) );
  NAND2_X2 U9630 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  NAND2_X2 U9631 ( .A1(n7508), .A2(n7507), .ZN(n7748) );
  INV_X4 U9632 ( .A(n7507), .ZN(n7510) );
  INV_X4 U9633 ( .A(n7508), .ZN(n7509) );
  NAND2_X2 U9634 ( .A1(n7510), .A2(n7509), .ZN(n7747) );
  NAND2_X2 U9635 ( .A1(a[16]), .A2(b[14]), .ZN(n7745) );
  XNOR2_X2 U9636 ( .A(n7511), .B(n7745), .ZN(n7751) );
  INV_X4 U9637 ( .A(n7513), .ZN(n7515) );
  OAI21_X4 U9638 ( .B1(n7342), .B2(n7515), .A(n7514), .ZN(n7752) );
  XNOR2_X2 U9639 ( .A(n7751), .B(n7752), .ZN(n7590) );
  INV_X4 U9640 ( .A(n7517), .ZN(n7519) );
  NAND2_X2 U9641 ( .A1(n7523), .A2(n3789), .ZN(n7760) );
  NAND2_X2 U9642 ( .A1(a[14]), .A2(b[16]), .ZN(n7758) );
  XNOR2_X2 U9643 ( .A(n7524), .B(n7758), .ZN(n7764) );
  INV_X4 U9644 ( .A(n7526), .ZN(n7528) );
  XNOR2_X2 U9645 ( .A(n7764), .B(n7765), .ZN(n7586) );
  NAND2_X2 U9646 ( .A1(a[13]), .A2(b[17]), .ZN(n7585) );
  XNOR2_X2 U9647 ( .A(n7586), .B(n7585), .ZN(n7534) );
  NAND2_X2 U9648 ( .A1(n7534), .A2(n7533), .ZN(n7773) );
  INV_X4 U9649 ( .A(n7533), .ZN(n7536) );
  INV_X4 U9650 ( .A(n7534), .ZN(n7535) );
  NAND2_X2 U9651 ( .A1(n7536), .A2(n7535), .ZN(n7772) );
  NAND2_X2 U9652 ( .A1(a[12]), .A2(b[18]), .ZN(n7770) );
  XNOR2_X2 U9653 ( .A(n7537), .B(n7770), .ZN(n7776) );
  XNOR2_X2 U9654 ( .A(n7776), .B(n3900), .ZN(n7583) );
  OAI21_X4 U9655 ( .B1(n7545), .B2(n3807), .A(n7543), .ZN(n7546) );
  NAND2_X2 U9656 ( .A1(n7547), .A2(n7546), .ZN(n7786) );
  INV_X4 U9657 ( .A(n7546), .ZN(n7548) );
  NAND2_X2 U9658 ( .A1(n7548), .A2(n3879), .ZN(n7785) );
  XNOR2_X2 U9659 ( .A(n7549), .B(n7783), .ZN(n7789) );
  XNOR2_X2 U9660 ( .A(n7789), .B(n7790), .ZN(n7579) );
  NAND2_X2 U9661 ( .A1(a[9]), .A2(b[21]), .ZN(n7578) );
  XNOR2_X2 U9662 ( .A(n7579), .B(n7578), .ZN(n7557) );
  NAND2_X2 U9663 ( .A1(n7556), .A2(n7557), .ZN(n7581) );
  INV_X4 U9664 ( .A(n7556), .ZN(n7559) );
  INV_X4 U9665 ( .A(n7557), .ZN(n7558) );
  NAND2_X2 U9666 ( .A1(n7559), .A2(n7558), .ZN(n7574) );
  NAND2_X2 U9667 ( .A1(n7581), .A2(n7574), .ZN(n7560) );
  XNOR2_X2 U9668 ( .A(net212146), .B(n7560), .ZN(n7562) );
  NAND2_X2 U9669 ( .A1(a[7]), .A2(b[23]), .ZN(n7575) );
  NAND2_X2 U9670 ( .A1(b[22]), .A2(a[8]), .ZN(n7795) );
  XNOR2_X2 U9671 ( .A(n7575), .B(n7795), .ZN(n7561) );
  XNOR2_X2 U9672 ( .A(n7562), .B(n7561), .ZN(n7563) );
  NAND2_X2 U9673 ( .A1(n7563), .A2(net212451), .ZN(net212137) );
  INV_X4 U9674 ( .A(n7563), .ZN(n7564) );
  NAND2_X2 U9675 ( .A1(net212448), .A2(n7564), .ZN(net212138) );
  NAND2_X2 U9676 ( .A1(b[24]), .A2(a[6]), .ZN(net212140) );
  XNOR2_X2 U9677 ( .A(net212447), .B(net212140), .ZN(n7801) );
  XNOR2_X2 U9678 ( .A(n7565), .B(n7801), .ZN(n7567) );
  NAND2_X2 U9679 ( .A1(n7566), .A2(n7567), .ZN(net212126) );
  INV_X4 U9680 ( .A(n7566), .ZN(n7570) );
  INV_X4 U9681 ( .A(n7567), .ZN(n7569) );
  NAND2_X2 U9682 ( .A1(net219055), .A2(b[26]), .ZN(net212128) );
  NAND2_X2 U9683 ( .A1(a[3]), .A2(b[27]), .ZN(net212393) );
  XNOR2_X2 U9684 ( .A(net212433), .B(net212128), .ZN(net212121) );
  INV_X4 U9685 ( .A(net212121), .ZN(net212394) );
  NAND2_X2 U9686 ( .A1(n7570), .A2(n7569), .ZN(net212125) );
  INV_X4 U9687 ( .A(net212125), .ZN(net212383) );
  NOR2_X2 U9688 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  NOR2_X4 U9689 ( .A1(net212383), .A2(n7573), .ZN(net212129) );
  NAND2_X2 U9690 ( .A1(n7581), .A2(n7574), .ZN(n7796) );
  XNOR2_X2 U9691 ( .A(n7796), .B(n7795), .ZN(net212381) );
  INV_X4 U9692 ( .A(net212381), .ZN(net212145) );
  NOR2_X4 U9693 ( .A1(net212377), .A2(n7577), .ZN(net212141) );
  INV_X4 U9694 ( .A(n7578), .ZN(n7580) );
  NAND2_X2 U9695 ( .A1(n7582), .A2(n7581), .ZN(n7794) );
  NAND2_X2 U9696 ( .A1(n7584), .A2(n7786), .ZN(n7782) );
  INV_X4 U9697 ( .A(n7585), .ZN(n7587) );
  NAND2_X2 U9698 ( .A1(n7591), .A2(n7590), .ZN(n7592) );
  NAND2_X2 U9699 ( .A1(n7592), .A2(n7761), .ZN(n7757) );
  INV_X4 U9700 ( .A(n7593), .ZN(n7596) );
  XNOR2_X2 U9701 ( .A(n7594), .B(n7599), .ZN(n7595) );
  NAND2_X2 U9702 ( .A1(n7596), .A2(n7595), .ZN(n7597) );
  NAND2_X2 U9703 ( .A1(n7597), .A2(n7748), .ZN(n7744) );
  NAND2_X2 U9704 ( .A1(n7599), .A2(n7598), .ZN(n7742) );
  INV_X4 U9705 ( .A(n7600), .ZN(n7603) );
  XNOR2_X2 U9706 ( .A(n7730), .B(n7601), .ZN(n7602) );
  NAND2_X2 U9707 ( .A1(n7603), .A2(n7602), .ZN(n7605) );
  NAND2_X2 U9708 ( .A1(n7605), .A2(n7604), .ZN(n7734) );
  INV_X4 U9709 ( .A(n7606), .ZN(n7608) );
  NOR2_X4 U9710 ( .A1(n7608), .A2(n7607), .ZN(n7728) );
  INV_X4 U9711 ( .A(n7612), .ZN(n7614) );
  NOR2_X4 U9712 ( .A1(n7614), .A2(n7613), .ZN(n7722) );
  INV_X4 U9713 ( .A(n7615), .ZN(n7616) );
  INV_X4 U9714 ( .A(n7619), .ZN(n7621) );
  NOR2_X4 U9715 ( .A1(n7621), .A2(n7620), .ZN(n7716) );
  INV_X4 U9716 ( .A(n7622), .ZN(n7626) );
  INV_X4 U9717 ( .A(n7623), .ZN(n7625) );
  INV_X4 U9718 ( .A(n7627), .ZN(n7710) );
  INV_X4 U9719 ( .A(n7628), .ZN(n7629) );
  INV_X4 U9720 ( .A(n7632), .ZN(n7636) );
  INV_X4 U9721 ( .A(n7633), .ZN(n7635) );
  OAI21_X4 U9722 ( .B1(n7636), .B2(n7635), .A(n7634), .ZN(n7706) );
  NAND2_X2 U9723 ( .A1(n7638), .A2(n7637), .ZN(n7704) );
  NAND2_X2 U9724 ( .A1(a[19]), .A2(b[12]), .ZN(n7640) );
  NAND2_X2 U9725 ( .A1(a[13]), .A2(b[18]), .ZN(n7639) );
  XOR2_X2 U9726 ( .A(n7640), .B(n7639), .Z(n7644) );
  NAND2_X2 U9727 ( .A1(a[22]), .A2(b[9]), .ZN(n7642) );
  NAND2_X2 U9728 ( .A1(a[10]), .A2(b[21]), .ZN(n7641) );
  XNOR2_X2 U9729 ( .A(n7642), .B(n7641), .ZN(n7643) );
  XNOR2_X2 U9730 ( .A(n7644), .B(n7643), .ZN(n7652) );
  NAND2_X2 U9731 ( .A1(a[21]), .A2(b[10]), .ZN(n7646) );
  NAND2_X2 U9732 ( .A1(a[12]), .A2(b[19]), .ZN(n7645) );
  XOR2_X2 U9733 ( .A(n7646), .B(n7645), .Z(n7650) );
  NAND2_X2 U9734 ( .A1(a[24]), .A2(b[7]), .ZN(n7648) );
  NAND2_X2 U9735 ( .A1(a[11]), .A2(b[20]), .ZN(n7647) );
  XNOR2_X2 U9736 ( .A(n7648), .B(n7647), .ZN(n7649) );
  XNOR2_X2 U9737 ( .A(n7650), .B(n7649), .ZN(n7651) );
  XNOR2_X2 U9738 ( .A(n7652), .B(n7651), .ZN(n7666) );
  NAND2_X2 U9739 ( .A1(a[20]), .A2(b[11]), .ZN(n7654) );
  NAND2_X2 U9740 ( .A1(a[17]), .A2(b[14]), .ZN(n7653) );
  XNOR2_X2 U9741 ( .A(n7654), .B(n7653), .ZN(n7658) );
  NAND2_X2 U9742 ( .A1(a[14]), .A2(b[17]), .ZN(n7656) );
  NAND2_X2 U9743 ( .A1(a[16]), .A2(b[15]), .ZN(n7655) );
  XNOR2_X2 U9744 ( .A(n7656), .B(n7655), .ZN(n7657) );
  XNOR2_X2 U9745 ( .A(n7658), .B(n7657), .ZN(n7664) );
  NAND2_X2 U9746 ( .A1(b[13]), .A2(a[18]), .ZN(n7660) );
  NAND2_X2 U9747 ( .A1(a[15]), .A2(b[16]), .ZN(n7659) );
  XNOR2_X2 U9748 ( .A(n7660), .B(n7659), .ZN(n7662) );
  NAND2_X2 U9749 ( .A1(a[29]), .A2(net218550), .ZN(n7661) );
  XNOR2_X2 U9750 ( .A(n7662), .B(n7661), .ZN(n7663) );
  XNOR2_X2 U9751 ( .A(n7664), .B(n7663), .ZN(n7665) );
  XNOR2_X2 U9752 ( .A(n7666), .B(n7665), .ZN(n7672) );
  NOR2_X4 U9753 ( .A1(net218624), .A2(net212284), .ZN(n7667) );
  MUX2_X2 U9754 ( .A(n7668), .B(n7667), .S(a[30]), .Z(n7670) );
  NAND2_X2 U9755 ( .A1(n7670), .A2(n7669), .ZN(n7671) );
  XNOR2_X2 U9756 ( .A(n7672), .B(n7671), .ZN(n7702) );
  NAND2_X2 U9757 ( .A1(a[8]), .A2(b[23]), .ZN(n7674) );
  NAND2_X2 U9758 ( .A1(a[25]), .A2(b[6]), .ZN(n7673) );
  XOR2_X2 U9759 ( .A(n7674), .B(n7673), .Z(n7678) );
  NAND2_X2 U9760 ( .A1(b[25]), .A2(a[6]), .ZN(n7676) );
  NAND2_X2 U9761 ( .A1(a[23]), .A2(b[8]), .ZN(n7675) );
  XNOR2_X2 U9762 ( .A(n7676), .B(n7675), .ZN(n7677) );
  XNOR2_X2 U9763 ( .A(n7678), .B(n7677), .ZN(n7686) );
  NAND2_X2 U9764 ( .A1(a[5]), .A2(b[26]), .ZN(n7680) );
  NAND2_X2 U9765 ( .A1(b[24]), .A2(a[7]), .ZN(n7679) );
  XNOR2_X2 U9766 ( .A(n7680), .B(n7679), .ZN(n7684) );
  NAND2_X2 U9767 ( .A1(a[26]), .A2(b[5]), .ZN(n7682) );
  NAND2_X2 U9768 ( .A1(b[22]), .A2(a[9]), .ZN(n7681) );
  XNOR2_X2 U9769 ( .A(n7682), .B(n7681), .ZN(n7683) );
  XNOR2_X2 U9770 ( .A(n7684), .B(n7683), .ZN(n7685) );
  XNOR2_X2 U9771 ( .A(n7686), .B(n7685), .ZN(n7700) );
  NAND2_X2 U9772 ( .A1(b[29]), .A2(a[2]), .ZN(n7687) );
  XOR2_X2 U9773 ( .A(n7688), .B(n7687), .Z(n7692) );
  NAND2_X2 U9774 ( .A1(a[27]), .A2(b[4]), .ZN(n7690) );
  NAND2_X2 U9775 ( .A1(b[28]), .A2(a[3]), .ZN(n7689) );
  XNOR2_X2 U9776 ( .A(n7690), .B(n7689), .ZN(n7691) );
  XNOR2_X2 U9777 ( .A(n7692), .B(n7691), .ZN(n7698) );
  NAND2_X2 U9778 ( .A1(a[28]), .A2(net218540), .ZN(n7694) );
  XNOR2_X2 U9779 ( .A(n7694), .B(n7693), .ZN(n7696) );
  XNOR2_X2 U9780 ( .A(n7696), .B(n7695), .ZN(n7697) );
  XNOR2_X2 U9781 ( .A(n7698), .B(n7697), .ZN(n7699) );
  XNOR2_X2 U9782 ( .A(n7700), .B(n7699), .ZN(n7701) );
  XNOR2_X2 U9783 ( .A(n7702), .B(n7701), .ZN(n7703) );
  XNOR2_X2 U9784 ( .A(n7704), .B(n7703), .ZN(n7705) );
  XNOR2_X2 U9785 ( .A(n7706), .B(n7705), .ZN(n7707) );
  XNOR2_X2 U9786 ( .A(n7708), .B(n7707), .ZN(n7709) );
  XNOR2_X2 U9787 ( .A(n7710), .B(n7709), .ZN(n7712) );
  XNOR2_X2 U9788 ( .A(n7712), .B(n7711), .ZN(n7713) );
  XNOR2_X2 U9789 ( .A(n7714), .B(n7713), .ZN(n7715) );
  XNOR2_X2 U9790 ( .A(n7716), .B(n7715), .ZN(n7717) );
  XNOR2_X2 U9791 ( .A(n7718), .B(n7717), .ZN(n7719) );
  XNOR2_X2 U9792 ( .A(n7720), .B(n7719), .ZN(n7721) );
  XNOR2_X2 U9793 ( .A(n7722), .B(n7721), .ZN(n7724) );
  XNOR2_X2 U9794 ( .A(n7724), .B(n7723), .ZN(n7725) );
  XNOR2_X2 U9795 ( .A(n7726), .B(n7725), .ZN(n7727) );
  XNOR2_X2 U9796 ( .A(n7728), .B(n7727), .ZN(n7732) );
  NOR2_X4 U9797 ( .A1(n7730), .A2(n7729), .ZN(n7731) );
  XNOR2_X2 U9798 ( .A(n7732), .B(n7731), .ZN(n7733) );
  XNOR2_X2 U9799 ( .A(n7734), .B(n7733), .ZN(n7740) );
  INV_X4 U9800 ( .A(n7735), .ZN(n7738) );
  INV_X4 U9801 ( .A(n7736), .ZN(n7737) );
  NAND2_X2 U9802 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  XNOR2_X2 U9803 ( .A(n7740), .B(n7739), .ZN(n7741) );
  XNOR2_X2 U9804 ( .A(n7742), .B(n7741), .ZN(n7743) );
  XNOR2_X2 U9805 ( .A(n7744), .B(n7743), .ZN(n7750) );
  INV_X4 U9806 ( .A(n7745), .ZN(n7746) );
  NAND3_X2 U9807 ( .A1(n7748), .A2(n7747), .A3(n7746), .ZN(n7749) );
  XNOR2_X2 U9808 ( .A(n7750), .B(n7749), .ZN(n7755) );
  INV_X4 U9809 ( .A(n7751), .ZN(n7753) );
  NAND2_X2 U9810 ( .A1(n7753), .A2(n7752), .ZN(n7754) );
  XNOR2_X2 U9811 ( .A(n7755), .B(n7754), .ZN(n7756) );
  XNOR2_X2 U9812 ( .A(n7757), .B(n7756), .ZN(n7763) );
  INV_X4 U9813 ( .A(n7758), .ZN(n7759) );
  NAND3_X2 U9814 ( .A1(n7761), .A2(n7760), .A3(n7759), .ZN(n7762) );
  XNOR2_X2 U9815 ( .A(n7763), .B(n7762), .ZN(n7767) );
  XNOR2_X2 U9816 ( .A(n7767), .B(n7766), .ZN(n7768) );
  XNOR2_X2 U9817 ( .A(n7769), .B(n7768), .ZN(n7775) );
  INV_X4 U9818 ( .A(n7770), .ZN(n7771) );
  XNOR2_X2 U9819 ( .A(n7775), .B(n7774), .ZN(n7780) );
  INV_X4 U9820 ( .A(n3919), .ZN(n7778) );
  NAND2_X2 U9821 ( .A1(n7778), .A2(n3900), .ZN(n7779) );
  XNOR2_X2 U9822 ( .A(n7780), .B(n7779), .ZN(n7781) );
  XNOR2_X2 U9823 ( .A(n7782), .B(n7781), .ZN(n7788) );
  INV_X4 U9824 ( .A(n7783), .ZN(n7784) );
  XNOR2_X2 U9825 ( .A(n7788), .B(n7787), .ZN(n7792) );
  NAND2_X2 U9826 ( .A1(n3896), .A2(n7790), .ZN(n7791) );
  XNOR2_X2 U9827 ( .A(n7792), .B(n7791), .ZN(n7793) );
  XNOR2_X2 U9828 ( .A(n7794), .B(n7793), .ZN(n7800) );
  INV_X4 U9829 ( .A(n7795), .ZN(n7798) );
  INV_X4 U9830 ( .A(n7796), .ZN(n7797) );
  NAND2_X2 U9831 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  XNOR2_X2 U9832 ( .A(n7800), .B(n7799), .ZN(net212143) );
  AOI21_X2 U9833 ( .B1(net218655), .B2(net218610), .A(net212023), .ZN(
        net212102) );
  NAND2_X2 U9834 ( .A1(net212093), .A2(net212094), .ZN(net212092) );
  NAND2_X2 U9835 ( .A1(n7803), .A2(n7802), .ZN(n7810) );
  NAND2_X2 U9836 ( .A1(n7805), .A2(n7804), .ZN(n7809) );
  NAND2_X2 U9837 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND3_X2 U9838 ( .A1(n7810), .A2(n7809), .A3(n7808), .ZN(n7812) );
  MUX2_X2 U9839 ( .A(n7812), .B(n7811), .S(b[4]), .Z(n7823) );
  INV_X4 U9840 ( .A(n7813), .ZN(n7814) );
  NOR2_X4 U9841 ( .A1(n7815), .A2(n7814), .ZN(n7820) );
  MUX2_X2 U9842 ( .A(n7817), .B(n7816), .S(net218558), .Z(n7819) );
  OAI21_X4 U9843 ( .B1(n7823), .B2(n7822), .A(n7821), .ZN(n7824) );
  INV_X4 U9844 ( .A(n7824), .ZN(n7892) );
  NOR2_X4 U9845 ( .A1(n7825), .A2(net218640), .ZN(n7827) );
  NOR2_X4 U9846 ( .A1(n7827), .A2(n7826), .ZN(n7833) );
  INV_X4 U9847 ( .A(n7828), .ZN(n7830) );
  AOI22_X2 U9848 ( .A1(n7856), .A2(n7831), .B1(n7830), .B2(n7829), .ZN(n7832)
         );
  NAND3_X2 U9849 ( .A1(n7833), .A2(n7832), .A3(net212061), .ZN(n7891) );
  NOR4_X2 U9850 ( .A1(result[2]), .A2(n7892), .A3(result[1]), .A4(n7891), .ZN(
        n7835) );
  INV_X4 U9851 ( .A(result[3]), .ZN(n7834) );
  NAND2_X2 U9852 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  NOR2_X4 U9853 ( .A1(result[8]), .A2(n3356), .ZN(n7838) );
  INV_X4 U9854 ( .A(result[0]), .ZN(n7837) );
  NAND2_X2 U9855 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  NOR2_X4 U9856 ( .A1(result[11]), .A2(n3358), .ZN(n7845) );
  XNOR2_X2 U9857 ( .A(n4002), .B(b[30]), .ZN(n7848) );
  XNOR2_X2 U9858 ( .A(n7848), .B(n7889), .ZN(n7847) );
  INV_X4 U9859 ( .A(a[29]), .ZN(n7842) );
  OAI22_X2 U9860 ( .A1(n7843), .A2(n7842), .B1(n7841), .B2(n7840), .ZN(n7850)
         );
  XNOR2_X2 U9861 ( .A(n7847), .B(n7850), .ZN(n7844) );
  NAND2_X2 U9862 ( .A1(n7844), .A2(n3990), .ZN(n7893) );
  NAND2_X2 U9863 ( .A1(n7845), .A2(n7893), .ZN(n7846) );
  NOR2_X4 U9864 ( .A1(result[12]), .A2(n7846), .ZN(n7886) );
  INV_X4 U9865 ( .A(n7847), .ZN(n7851) );
  XNOR2_X2 U9866 ( .A(n4002), .B(net211993), .ZN(n7852) );
  XNOR2_X2 U9867 ( .A(n7853), .B(n7852), .ZN(n7854) );
  NAND2_X2 U9868 ( .A1(n7854), .A2(n3990), .ZN(n7885) );
  NAND2_X2 U9869 ( .A1(n7856), .A2(n3998), .ZN(n7860) );
  NOR2_X4 U9870 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  NAND3_X2 U9871 ( .A1(n7860), .A2(net218610), .A3(n7859), .ZN(n7861) );
  NAND2_X2 U9872 ( .A1(a[31]), .A2(n7861), .ZN(n7884) );
  NAND2_X2 U9873 ( .A1(n7863), .A2(n7862), .ZN(n7868) );
  NAND2_X2 U9874 ( .A1(n7865), .A2(n7864), .ZN(n7867) );
  INV_X4 U9875 ( .A(net212010), .ZN(net212008) );
  INV_X4 U9876 ( .A(net212007), .ZN(net212005) );
  NOR3_X4 U9877 ( .A1(n7875), .A2(n7874), .A3(n7873), .ZN(n7877) );
  MUX2_X2 U9878 ( .A(n7877), .B(n7876), .S(b[4]), .Z(n7879) );
  AOI21_X2 U9879 ( .B1(n7880), .B2(n7879), .A(n7878), .ZN(n7882) );
  NOR2_X4 U9880 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  NAND2_X2 U9881 ( .A1(n7886), .A2(n3355), .ZN(n7887) );
endmodule

